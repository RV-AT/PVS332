module prv332sv0 ( gnd, vdd, clk, rst, timer_int, soft_int, ext_int, hready, hresp, hreset_n, hrdata, haddr, hwrite, hsize, hburst, hprot, htrans, hmastlock, hwdata);

input gnd, vdd;
input clk;
input rst;
input timer_int;
input soft_int;
input ext_int;
input hready;
input hresp;
input hreset_n;
output hwrite;
output hmastlock;
input [31:0] hrdata;
output [33:0] haddr;
output [1:0] hsize;
output [2:0] hburst;
output [3:0] hprot;
output [1:0] htrans;
output [31:0] hwdata;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf11) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf10) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf9) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
	BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
	BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
	BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3), .Y(_7303__bF_buf3_bF_buf3) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3), .Y(_7303__bF_buf3_bF_buf2) );
	BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3), .Y(_7303__bF_buf3_bF_buf1) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3), .Y(_7303__bF_buf3_bF_buf0) );
	BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4), .Y(_7303__bF_buf4_bF_buf3) );
	BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4), .Y(_7303__bF_buf4_bF_buf2) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4), .Y(_7303__bF_buf4_bF_buf1) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4), .Y(_7303__bF_buf4_bF_buf0) );
	BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5), .Y(_7303__bF_buf5_bF_buf3) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5), .Y(_7303__bF_buf5_bF_buf2) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5), .Y(_7303__bF_buf5_bF_buf1) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5), .Y(_7303__bF_buf5_bF_buf0) );
	BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6), .Y(_7303__bF_buf6_bF_buf3) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6), .Y(_7303__bF_buf6_bF_buf2) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6), .Y(_7303__bF_buf6_bF_buf1) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6), .Y(_7303__bF_buf6_bF_buf0) );
	BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7), .Y(_7303__bF_buf7_bF_buf3) );
	BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7), .Y(_7303__bF_buf7_bF_buf2) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7), .Y(_7303__bF_buf7_bF_buf1) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7), .Y(_7303__bF_buf7_bF_buf0) );
	BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8), .Y(_7303__bF_buf8_bF_buf3) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8), .Y(_7303__bF_buf8_bF_buf2) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8), .Y(_7303__bF_buf8_bF_buf1) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8), .Y(_7303__bF_buf8_bF_buf0) );
	BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9), .Y(_7303__bF_buf9_bF_buf3) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9), .Y(_7303__bF_buf9_bF_buf2) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9), .Y(_7303__bF_buf9_bF_buf1) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9), .Y(_7303__bF_buf9_bF_buf0) );
	BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10), .Y(_7304__bF_buf10_bF_buf3) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10), .Y(_7304__bF_buf10_bF_buf2) );
	BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10), .Y(_7304__bF_buf10_bF_buf1) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10), .Y(_7304__bF_buf10_bF_buf0) );
	BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11), .Y(_7304__bF_buf11_bF_buf3) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11), .Y(_7304__bF_buf11_bF_buf2) );
	BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11), .Y(_7304__bF_buf11_bF_buf1) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11), .Y(_7304__bF_buf11_bF_buf0) );
	BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12), .Y(_7304__bF_buf12_bF_buf3) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12), .Y(_7304__bF_buf12_bF_buf2) );
	BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12), .Y(_7304__bF_buf12_bF_buf1) );
	BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12), .Y(_7304__bF_buf12_bF_buf0) );
	BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13), .Y(_7304__bF_buf13_bF_buf3) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13), .Y(_7304__bF_buf13_bF_buf2) );
	BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13), .Y(_7304__bF_buf13_bF_buf1) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13), .Y(_7304__bF_buf13_bF_buf0) );
	BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14), .Y(_7304__bF_buf14_bF_buf3) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14), .Y(_7304__bF_buf14_bF_buf2) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14), .Y(_7304__bF_buf14_bF_buf1) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14), .Y(_7304__bF_buf14_bF_buf0) );
	BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6), .Y(_7304__bF_buf6_bF_buf3) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6), .Y(_7304__bF_buf6_bF_buf2) );
	BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6), .Y(_7304__bF_buf6_bF_buf1) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6), .Y(_7304__bF_buf6_bF_buf0) );
	BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7), .Y(_7304__bF_buf7_bF_buf3) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7), .Y(_7304__bF_buf7_bF_buf2) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7), .Y(_7304__bF_buf7_bF_buf1) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7), .Y(_7304__bF_buf7_bF_buf0) );
	BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8), .Y(_7304__bF_buf8_bF_buf3) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8), .Y(_7304__bF_buf8_bF_buf2) );
	BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8), .Y(_7304__bF_buf8_bF_buf1) );
	BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8), .Y(_7304__bF_buf8_bF_buf0) );
	BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9), .Y(_7304__bF_buf9_bF_buf3) );
	BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9), .Y(_7304__bF_buf9_bF_buf2) );
	BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9), .Y(_7304__bF_buf9_bF_buf1) );
	BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9), .Y(_7304__bF_buf9_bF_buf0) );
	BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf5) );
	BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf4) );
	BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf3) );
	BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf2) );
	BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf1) );
	BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6879__hier0_bF_buf0) );
	BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10), .Y(_7303__bF_buf10_bF_buf3) );
	BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10), .Y(_7303__bF_buf10_bF_buf2) );
	BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10), .Y(_7303__bF_buf10_bF_buf1) );
	BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10), .Y(_7303__bF_buf10_bF_buf0) );
	BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11), .Y(_7303__bF_buf11_bF_buf3) );
	BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11), .Y(_7303__bF_buf11_bF_buf2) );
	BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11), .Y(_7303__bF_buf11_bF_buf1) );
	BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11), .Y(_7303__bF_buf11_bF_buf0) );
	BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12), .Y(_7303__bF_buf12_bF_buf3) );
	BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12), .Y(_7303__bF_buf12_bF_buf2) );
	BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12), .Y(_7303__bF_buf12_bF_buf1) );
	BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12), .Y(_7303__bF_buf12_bF_buf0) );
	BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13), .Y(_7303__bF_buf13_bF_buf3) );
	BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13), .Y(_7303__bF_buf13_bF_buf2) );
	BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13), .Y(_7303__bF_buf13_bF_buf1) );
	BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13), .Y(_7303__bF_buf13_bF_buf0) );
	BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14), .Y(_7303__bF_buf14_bF_buf3) );
	BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14), .Y(_7303__bF_buf14_bF_buf2) );
	BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14), .Y(_7303__bF_buf14_bF_buf1) );
	BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14), .Y(_7303__bF_buf14_bF_buf0) );
	BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf7) );
	BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf6) );
	BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf5) );
	BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf4) );
	BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf3) );
	BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf2) );
	BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf1) );
	BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_hier0_bF_buf0) );
	BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7434__bF_buf4) );
	BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7434__bF_buf3) );
	BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7434__bF_buf2) );
	BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7434__bF_buf1) );
	BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7434__bF_buf0) );
	BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_32__bF_buf3) );
	BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_32__bF_buf2) );
	BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_32__bF_buf1) );
	BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_32__bF_buf0) );
	BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .Y(_6292__bF_buf4) );
	BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .Y(_6292__bF_buf3) );
	BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .Y(_6292__bF_buf2) );
	BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .Y(_6292__bF_buf1) );
	BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .Y(_6292__bF_buf0) );
	BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf10) );
	BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf9) );
	BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf8) );
	BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf7) );
	BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf6) );
	BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf5) );
	BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf4) );
	BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf3) );
	BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf2) );
	BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf1) );
	BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .Y(_6160__bF_buf0) );
	BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .Y(_14545__bF_buf3) );
	BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .Y(_14545__bF_buf2) );
	BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .Y(_14545__bF_buf1) );
	BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .Y(_14545__bF_buf0) );
	BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2499__bF_buf4) );
	BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2499__bF_buf3) );
	BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2499__bF_buf2) );
	BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2499__bF_buf1) );
	BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2499__bF_buf0) );
	BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_13776_), .Y(_13776__bF_buf3) );
	BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_13776_), .Y(_13776__bF_buf2) );
	BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_13776_), .Y(_13776__bF_buf1) );
	BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_13776_), .Y(_13776__bF_buf0) );
	BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .Y(_6931__bF_buf3) );
	BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .Y(_6931__bF_buf2) );
	BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .Y(_6931__bF_buf1) );
	BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .Y(_6931__bF_buf0) );
	BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf6) );
	BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf5) );
	BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf4) );
	BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf3) );
	BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf2) );
	BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf1) );
	BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .Y(_13415__bF_buf0) );
	BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1068__bF_buf4) );
	BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1068__bF_buf3) );
	BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1068__bF_buf2) );
	BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1068__bF_buf1) );
	BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1068__bF_buf0) );
	BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf5) );
	BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf4) );
	BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf3) );
	BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf2) );
	BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf1) );
	BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .Y(_4893__bF_buf0) );
	BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .Y(_13470__bF_buf4) );
	BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .Y(_13470__bF_buf3) );
	BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .Y(_13470__bF_buf2) );
	BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .Y(_13470__bF_buf1) );
	BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .Y(_13470__bF_buf0) );
	BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf5) );
	BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf4) );
	BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf3) );
	BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf2) );
	BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf1) );
	BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .Y(_8328__bF_buf0) );
	BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2994__bF_buf4) );
	BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2994__bF_buf3) );
	BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2994__bF_buf2) );
	BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2994__bF_buf1) );
	BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2994__bF_buf0) );
	BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf5) );
	BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf4) );
	BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf3) );
	BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf2) );
	BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf1) );
	BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .Y(_8557__bF_buf0) );
	BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2862__bF_buf4) );
	BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2862__bF_buf3) );
	BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2862__bF_buf2) );
	BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2862__bF_buf1) );
	BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2862__bF_buf0) );
	BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2531__bF_buf4) );
	BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2531__bF_buf3) );
	BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2531__bF_buf2) );
	BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2531__bF_buf1) );
	BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2531__bF_buf0) );
	BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2501__bF_buf4) );
	BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2501__bF_buf3) );
	BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2501__bF_buf2) );
	BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2501__bF_buf1) );
	BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2501__bF_buf0) );
	BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .Y(_6459__bF_buf4) );
	BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .Y(_6459__bF_buf3) );
	BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .Y(_6459__bF_buf2) );
	BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .Y(_6459__bF_buf1) );
	BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .Y(_6459__bF_buf0) );
	BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf5) );
	BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf4) );
	BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf3) );
	BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf2) );
	BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf1) );
	BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .Y(_8684__bF_buf0) );
	BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf5) );
	BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf4) );
	BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf3) );
	BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf2) );
	BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf1) );
	BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_2730__bF_buf0) );
	BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .Y(_9020__bF_buf3) );
	BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .Y(_9020__bF_buf2) );
	BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .Y(_9020__bF_buf1) );
	BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .Y(_9020__bF_buf0) );
	BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf10) );
	BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf9) );
	BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf8) );
	BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf7) );
	BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf6) );
	BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf5) );
	BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf4) );
	BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf3) );
	BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf2) );
	BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf1) );
	BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .Y(_6026__bF_buf0) );
	BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf5) );
	BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf4) );
	BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf3) );
	BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf2) );
	BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf1) );
	BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .Y(_8281__bF_buf0) );
	BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf5) );
	BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf4) );
	BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf3) );
	BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf2) );
	BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf1) );
	BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .Y(_7584__bF_buf0) );
	BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf160) );
	BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf159) );
	BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf158) );
	BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf157) );
	BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf156) );
	BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf155) );
	BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf154) );
	BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf153) );
	BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf152) );
	BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf151) );
	BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf150) );
	BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf149) );
	BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf148) );
	BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf147) );
	BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf146) );
	BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf145) );
	BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf144) );
	BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf143) );
	BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf142) );
	BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf141) );
	BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf140) );
	BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf139) );
	BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf138) );
	BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf137) );
	BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf136) );
	BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf135) );
	BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf134) );
	BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf133) );
	BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf132) );
	BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf131) );
	BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf130) );
	BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf129) );
	BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf128) );
	BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf127) );
	BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf126) );
	BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf125) );
	BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf124) );
	BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf123) );
	BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf122) );
	BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf121) );
	BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf120) );
	BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf119) );
	BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf118) );
	BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf117) );
	BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf116) );
	BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf115) );
	BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf114) );
	BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf113) );
	BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf112) );
	BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf111) );
	BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf110) );
	BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf109) );
	BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf108) );
	BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf107) );
	BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf106) );
	BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf105) );
	BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf104) );
	BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf103) );
	BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf102) );
	BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf101) );
	BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf100) );
	BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf99) );
	BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf98) );
	BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf97) );
	BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf96) );
	BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf95) );
	BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf94) );
	BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf93) );
	BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf92) );
	BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf91) );
	BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf90) );
	BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf89) );
	BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf88) );
	BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf87) );
	BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf86) );
	BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf85) );
	BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf84) );
	BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf83) );
	BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf82) );
	BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf81) );
	BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf80) );
	BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf79) );
	BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf78) );
	BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf77) );
	BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf76) );
	BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf75) );
	BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf74) );
	BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf73) );
	BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf72) );
	BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf71) );
	BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf70) );
	BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf69) );
	BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf68) );
	BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf67) );
	BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf66) );
	BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf65) );
	BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf64) );
	BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf63) );
	BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf62) );
	BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf61) );
	BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf60) );
	BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf59) );
	BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf58) );
	BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57) );
	BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf56) );
	BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf55) );
	BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf54) );
	BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53) );
	BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf52) );
	BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf51) );
	BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf50) );
	BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf49) );
	BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf48) );
	BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf47) );
	BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf46) );
	BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf45) );
	BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf44) );
	BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf43) );
	BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf42) );
	BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf41) );
	BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf40) );
	BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf39) );
	BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf38) );
	BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf37) );
	BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf36) );
	BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf35) );
	BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf34) );
	BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf33) );
	BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf32) );
	BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf31) );
	BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf30) );
	BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf29) );
	BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf28) );
	BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf27) );
	BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf26) );
	BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25) );
	BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24) );
	BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23) );
	BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22) );
	BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf21) );
	BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20) );
	BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf19) );
	BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18) );
	BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17) );
	BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf16) );
	BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf15) );
	BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf14) );
	BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf13) );
	BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf12) );
	BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .Y(_7320__bF_buf3) );
	BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .Y(_7320__bF_buf2) );
	BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .Y(_7320__bF_buf1) );
	BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .Y(_7320__bF_buf0) );
	BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(_14334_), .Y(_14334__bF_buf4) );
	BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(_14334_), .Y(_14334__bF_buf3) );
	BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(_14334_), .Y(_14334__bF_buf2) );
	BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(_14334_), .Y(_14334__bF_buf1) );
	BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(_14334_), .Y(_14334__bF_buf0) );
	BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .Y(_4886__bF_buf3) );
	BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .Y(_4886__bF_buf2) );
	BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .Y(_4886__bF_buf1) );
	BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .Y(_4886__bF_buf0) );
	BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .Y(_2589__bF_buf4) );
	BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .Y(_2589__bF_buf3) );
	BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .Y(_2589__bF_buf2) );
	BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .Y(_2589__bF_buf1) );
	BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .Y(_2589__bF_buf0) );
	BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2529__bF_buf4) );
	BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2529__bF_buf3) );
	BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2529__bF_buf2) );
	BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2529__bF_buf1) );
	BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2529__bF_buf0) );
	BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf8) );
	BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf7) );
	BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf6) );
	BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf5) );
	BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf4) );
	BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf3) );
	BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf2) );
	BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf1) );
	BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2487__bF_buf0) );
	BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .Y(_13463__bF_buf4) );
	BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .Y(_13463__bF_buf3) );
	BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .Y(_13463__bF_buf2) );
	BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .Y(_13463__bF_buf1) );
	BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .Y(_13463__bF_buf0) );
	BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf7) );
	BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf6) );
	BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf5) );
	BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf4) );
	BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf3) );
	BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf2) );
	BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf1) );
	BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .Y(_13391__bF_buf0) );
	BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf11) );
	BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf10) );
	BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf9) );
	BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf8) );
	BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf7) );
	BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf6) );
	BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf5) );
	BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf4) );
	BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf3) );
	BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf2) );
	BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf1) );
	BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf0) );
	BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .Y(_9175__bF_buf4) );
	BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .Y(_9175__bF_buf3) );
	BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .Y(_9175__bF_buf2) );
	BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .Y(_9175__bF_buf1) );
	BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .Y(_9175__bF_buf0) );
	BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf5) );
	BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf4) );
	BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf3) );
	BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf2) );
	BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf1) );
	BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf0) );
	BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .Y(_12291__bF_buf3) );
	BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .Y(_12291__bF_buf2) );
	BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .Y(_12291__bF_buf1) );
	BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .Y(_12291__bF_buf0) );
	BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf6) );
	BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf5) );
	BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf4) );
	BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf3) );
	BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf2) );
	BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf1) );
	BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8117__bF_buf0) );
	BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .Y(_11402__bF_buf3) );
	BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .Y(_11402__bF_buf2) );
	BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .Y(_11402__bF_buf1) );
	BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .Y(_11402__bF_buf0) );
	BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_), .Y(biu_mmu_msu_0_bF_buf4) );
	BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_), .Y(biu_mmu_msu_0_bF_buf3) );
	BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_), .Y(biu_mmu_msu_0_bF_buf2) );
	BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_), .Y(biu_mmu_msu_0_bF_buf1) );
	BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_), .Y(biu_mmu_msu_0_bF_buf0) );
	BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(_8846_), .Y(_8846__bF_buf3) );
	BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(_8846_), .Y(_8846__bF_buf2) );
	BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(_8846_), .Y(_8846__bF_buf1) );
	BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(_8846_), .Y(_8846__bF_buf0) );
	BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .Y(_9110__bF_buf3) );
	BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .Y(_9110__bF_buf2) );
	BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .Y(_9110__bF_buf1) );
	BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .Y(_9110__bF_buf0) );
	BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf5) );
	BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf4) );
	BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf3) );
	BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf2) );
	BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf1) );
	BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .Y(_1220__bF_buf0) );
	BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf9) );
	BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf8) );
	BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf7) );
	BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf6) );
	BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf5) );
	BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf4) );
	BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf3) );
	BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf2) );
	BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf1) );
	BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .Y(_3117__bF_buf0) );
	BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_), .Y(biu_ins_25_bF_buf3) );
	BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_), .Y(biu_ins_25_bF_buf2) );
	BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_), .Y(biu_ins_25_bF_buf1) );
	BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_), .Y(biu_ins_25_bF_buf0) );
	BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_), .Y(addr_csr_27_bF_buf3) );
	BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_), .Y(addr_csr_27_bF_buf2) );
	BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_), .Y(addr_csr_27_bF_buf1) );
	BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_), .Y(addr_csr_27_bF_buf0) );
	BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf4) );
	BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf3) );
	BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf2) );
	BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf1) );
	BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf0) );
	BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .Y(_2517__bF_buf4) );
	BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .Y(_2517__bF_buf3) );
	BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .Y(_2517__bF_buf2) );
	BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .Y(_2517__bF_buf1) );
	BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .Y(_2517__bF_buf0) );
	BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(_14822_), .Y(_14822__bF_buf3) );
	BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(_14822_), .Y(_14822__bF_buf2) );
	BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_14822_), .Y(_14822__bF_buf1) );
	BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(_14822_), .Y(_14822__bF_buf0) );
	BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf6) );
	BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf5) );
	BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf4) );
	BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf3) );
	BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf2) );
	BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf1) );
	BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_), .Y(biu_ins_20_bF_buf0) );
	BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf5) );
	BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf4) );
	BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf3) );
	BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf2) );
	BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf1) );
	BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4911__bF_buf0) );
	BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_), .Y(csr_gpr_iu_csr_scause_31_bF_buf3) );
	BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_), .Y(csr_gpr_iu_csr_scause_31_bF_buf2) );
	BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_), .Y(csr_gpr_iu_csr_scause_31_bF_buf1) );
	BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_), .Y(csr_gpr_iu_csr_scause_31_bF_buf0) );
	BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .Y(_8165__bF_buf4) );
	BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .Y(_8165__bF_buf3) );
	BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .Y(_8165__bF_buf2) );
	BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .Y(_8165__bF_buf1) );
	BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .Y(_8165__bF_buf0) );
	BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(amoadd), .Y(amoadd_bF_buf3) );
	BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(amoadd), .Y(amoadd_bF_buf2) );
	BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(amoadd), .Y(amoadd_bF_buf1) );
	BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(amoadd), .Y(amoadd_bF_buf0) );
	BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf5) );
	BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf4) );
	BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf3) );
	BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf2) );
	BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf1) );
	BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8063__bF_buf0) );
	BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .Y(_7366__bF_buf3) );
	BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .Y(_7366__bF_buf2) );
	BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .Y(_7366__bF_buf1) );
	BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .Y(_7366__bF_buf0) );
	BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .Y(_6092__bF_buf4) );
	BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .Y(_6092__bF_buf3) );
	BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .Y(_6092__bF_buf2) );
	BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .Y(_6092__bF_buf1) );
	BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .Y(_6092__bF_buf0) );
	BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .Y(_6893__bF_buf4) );
	BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .Y(_6893__bF_buf3) );
	BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .Y(_6893__bF_buf2) );
	BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .Y(_6893__bF_buf1) );
	BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .Y(_6893__bF_buf0) );
	BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf15) );
	BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf14) );
	BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf13) );
	BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf12) );
	BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf11) );
	BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf10) );
	BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf9) );
	BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf8) );
	BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf7) );
	BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf6) );
	BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf5) );
	BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf4) );
	BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf3) );
	BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf2) );
	BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf1) );
	BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .Y(_4897__bF_buf0) );
	BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf7) );
	BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf6) );
	BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf5) );
	BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf4) );
	BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf3) );
	BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf2) );
	BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf1) );
	BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .Y(_3105__bF_buf0) );
	BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf5) );
	BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf4) );
	BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf3) );
	BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf2) );
	BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf1) );
	BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .Y(_6930__bF_buf0) );
	BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_), .Y(addr_csr_15_bF_buf3) );
	BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_), .Y(addr_csr_15_bF_buf2) );
	BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_), .Y(addr_csr_15_bF_buf1) );
	BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_), .Y(addr_csr_15_bF_buf0) );
	BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf5) );
	BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf4) );
	BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf3) );
	BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf2) );
	BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf1) );
	BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf0) );
	BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_14912__bF_buf4) );
	BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_14912__bF_buf3) );
	BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_14912__bF_buf2) );
	BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_14912__bF_buf1) );
	BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_14912__bF_buf0) );
	BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf5) );
	BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf4) );
	BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf3) );
	BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf2) );
	BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf1) );
	BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .Y(_8489__bF_buf0) );
	BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .Y(_2535__bF_buf4) );
	BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .Y(_2535__bF_buf3) );
	BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .Y(_2535__bF_buf2) );
	BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .Y(_2535__bF_buf1) );
	BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .Y(_2535__bF_buf0) );
	BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .Y(_2505__bF_buf4) );
	BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .Y(_2505__bF_buf3) );
	BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .Y(_2505__bF_buf2) );
	BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .Y(_2505__bF_buf1) );
	BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .Y(_2505__bF_buf0) );
	BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .Y(_2493__bF_buf4) );
	BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .Y(_2493__bF_buf3) );
	BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .Y(_2493__bF_buf2) );
	BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .Y(_2493__bF_buf1) );
	BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .Y(_2493__bF_buf0) );
	BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .Y(_3100__bF_buf3) );
	BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .Y(_3100__bF_buf2) );
	BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .Y(_3100__bF_buf1) );
	BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .Y(_3100__bF_buf0) );
	BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf6) );
	BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf5) );
	BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf4) );
	BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf3) );
	BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf2) );
	BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf1) );
	BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .Y(_8327__bF_buf0) );
	BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf5) );
	BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf4) );
	BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf3) );
	BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf2) );
	BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf1) );
	BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2993__bF_buf0) );
	BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .Y(_6259__bF_buf4) );
	BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .Y(_6259__bF_buf3) );
	BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .Y(_6259__bF_buf2) );
	BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .Y(_6259__bF_buf1) );
	BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .Y(_6259__bF_buf0) );
	BUFX4 BUFX4_619 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf12) );
	BUFX4 BUFX4_620 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf11) );
	BUFX4 BUFX4_621 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf10) );
	BUFX4 BUFX4_622 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf9) );
	BUFX4 BUFX4_623 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf8) );
	BUFX4 BUFX4_624 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf7) );
	BUFX4 BUFX4_625 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf6) );
	BUFX4 BUFX4_626 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf5) );
	BUFX4 BUFX4_627 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf4) );
	BUFX4 BUFX4_628 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf3) );
	BUFX4 BUFX4_629 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf2) );
	BUFX4 BUFX4_630 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf1) );
	BUFX4 BUFX4_631 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .Y(_2590__bF_buf0) );
	BUFX4 BUFX4_632 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .Y(_6759__bF_buf4) );
	BUFX4 BUFX4_633 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .Y(_6759__bF_buf3) );
	BUFX4 BUFX4_634 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .Y(_6759__bF_buf2) );
	BUFX4 BUFX4_635 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .Y(_6759__bF_buf1) );
	BUFX4 BUFX4_636 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .Y(_6759__bF_buf0) );
	BUFX4 BUFX4_637 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6326__bF_buf4) );
	BUFX4 BUFX4_638 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6326__bF_buf3) );
	BUFX4 BUFX4_639 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6326__bF_buf2) );
	BUFX4 BUFX4_640 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6326__bF_buf1) );
	BUFX4 BUFX4_641 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6326__bF_buf0) );
	BUFX4 BUFX4_642 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .Y(_6025__bF_buf4) );
	BUFX4 BUFX4_643 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .Y(_6025__bF_buf3) );
	BUFX4 BUFX4_644 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .Y(_6025__bF_buf2) );
	BUFX4 BUFX4_645 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .Y(_6025__bF_buf1) );
	BUFX4 BUFX4_646 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .Y(_6025__bF_buf0) );
	BUFX4 BUFX4_647 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf5) );
	BUFX4 BUFX4_648 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf4) );
	BUFX4 BUFX4_649 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf3) );
	BUFX4 BUFX4_650 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf2) );
	BUFX4 BUFX4_651 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf1) );
	BUFX4 BUFX4_652 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .Y(_8280__bF_buf0) );
	BUFX4 BUFX4_653 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .Y(_7583__bF_buf3) );
	BUFX4 BUFX4_654 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .Y(_7583__bF_buf2) );
	BUFX4 BUFX4_655 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .Y(_7583__bF_buf1) );
	BUFX4 BUFX4_656 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .Y(_7583__bF_buf0) );
	BUFX4 BUFX4_657 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .Y(_6525__bF_buf4) );
	BUFX4 BUFX4_658 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .Y(_6525__bF_buf3) );
	BUFX4 BUFX4_659 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .Y(_6525__bF_buf2) );
	BUFX4 BUFX4_660 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .Y(_6525__bF_buf1) );
	BUFX4 BUFX4_661 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .Y(_6525__bF_buf0) );
	BUFX4 BUFX4_662 ( .gnd(gnd), .vdd(vdd), .A(_6821_), .Y(_6821__bF_buf3) );
	BUFX4 BUFX4_663 ( .gnd(gnd), .vdd(vdd), .A(_6821_), .Y(_6821__bF_buf2) );
	BUFX4 BUFX4_664 ( .gnd(gnd), .vdd(vdd), .A(_6821_), .Y(_6821__bF_buf1) );
	BUFX4 BUFX4_665 ( .gnd(gnd), .vdd(vdd), .A(_6821_), .Y(_6821__bF_buf0) );
	BUFX4 BUFX4_666 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .Y(_12337__bF_buf3) );
	BUFX4 BUFX4_667 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .Y(_12337__bF_buf2) );
	BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .Y(_12337__bF_buf1) );
	BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .Y(_12337__bF_buf0) );
	BUFX4 BUFX4_668 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf7) );
	BUFX4 BUFX4_669 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf6) );
	BUFX4 BUFX4_670 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf5) );
	BUFX4 BUFX4_671 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf4) );
	BUFX4 BUFX4_672 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf3) );
	BUFX4 BUFX4_673 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf2) );
	BUFX4 BUFX4_674 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf1) );
	BUFX4 BUFX4_675 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .Y(_2588__bF_buf0) );
	BUFX4 BUFX4_676 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .Y(_9149__bF_buf4) );
	BUFX4 BUFX4_677 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .Y(_9149__bF_buf3) );
	BUFX4 BUFX4_678 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .Y(_9149__bF_buf2) );
	BUFX4 BUFX4_679 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .Y(_9149__bF_buf1) );
	BUFX4 BUFX4_680 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .Y(_9149__bF_buf0) );
	BUFX4 BUFX4_681 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf5) );
	BUFX4 BUFX4_682 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf4) );
	BUFX4 BUFX4_683 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf3) );
	BUFX4 BUFX4_684 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf2) );
	BUFX4 BUFX4_685 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf1) );
	BUFX4 BUFX4_686 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb), .Y(biu_ahb_rdy_ahb_bF_buf0) );
	BUFX4 BUFX4_687 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .Y(_13462__bF_buf3) );
	BUFX4 BUFX4_688 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .Y(_13462__bF_buf2) );
	BUFX4 BUFX4_689 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .Y(_13462__bF_buf1) );
	BUFX4 BUFX4_690 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .Y(_13462__bF_buf0) );
	BUFX4 BUFX4_691 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf6) );
	BUFX4 BUFX4_692 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf5) );
	BUFX4 BUFX4_693 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf4) );
	BUFX4 BUFX4_694 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf3) );
	BUFX4 BUFX4_695 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf2) );
	BUFX4 BUFX4_696 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf1) );
	BUFX4 BUFX4_697 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_), .Y(biu_ins_31_bF_buf0) );
	BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .Y(_9276__bF_buf3) );
	BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .Y(_9276__bF_buf2) );
	BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .Y(_9276__bF_buf1) );
	BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .Y(_9276__bF_buf0) );
	BUFX4 BUFX4_698 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2926__bF_buf4) );
	BUFX4 BUFX4_699 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2926__bF_buf3) );
	BUFX4 BUFX4_700 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2926__bF_buf2) );
	BUFX4 BUFX4_701 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2926__bF_buf1) );
	BUFX4 BUFX4_702 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2926__bF_buf0) );
	BUFX4 BUFX4_703 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf14) );
	BUFX4 BUFX4_704 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf13) );
	BUFX4 BUFX4_705 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf12) );
	BUFX4 BUFX4_706 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf11) );
	BUFX4 BUFX4_707 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf10) );
	BUFX4 BUFX4_708 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf9) );
	BUFX4 BUFX4_709 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf8) );
	BUFX4 BUFX4_710 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf7) );
	BUFX4 BUFX4_711 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf6) );
	BUFX4 BUFX4_712 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf5) );
	BUFX4 BUFX4_713 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf4) );
	BUFX4 BUFX4_714 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf3) );
	BUFX4 BUFX4_715 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf2) );
	BUFX4 BUFX4_716 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf1) );
	BUFX4 BUFX4_717 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .Y(_2625__bF_buf0) );
	BUFX4 BUFX4_718 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf10) );
	BUFX4 BUFX4_719 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf9) );
	BUFX4 BUFX4_720 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf8) );
	BUFX4 BUFX4_721 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf7) );
	BUFX4 BUFX4_722 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf6) );
	BUFX4 BUFX4_723 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf5) );
	BUFX4 BUFX4_724 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf4) );
	BUFX4 BUFX4_725 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf3) );
	BUFX4 BUFX4_726 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf2) );
	BUFX4 BUFX4_727 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf1) );
	BUFX4 BUFX4_728 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2553__bF_buf0) );
	BUFX4 BUFX4_729 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2523__bF_buf4) );
	BUFX4 BUFX4_730 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2523__bF_buf3) );
	BUFX4 BUFX4_731 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2523__bF_buf2) );
	BUFX4 BUFX4_732 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2523__bF_buf1) );
	BUFX4 BUFX4_733 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2523__bF_buf0) );
	BUFX4 BUFX4_734 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1224__bF_buf3) );
	BUFX4 BUFX4_735 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1224__bF_buf2) );
	BUFX4 BUFX4_736 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1224__bF_buf1) );
	BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1224__bF_buf0) );
	BUFX4 BUFX4_737 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .Y(_12290__bF_buf4) );
	BUFX4 BUFX4_738 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .Y(_12290__bF_buf3) );
	BUFX4 BUFX4_739 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .Y(_12290__bF_buf2) );
	BUFX4 BUFX4_740 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .Y(_12290__bF_buf1) );
	BUFX4 BUFX4_741 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .Y(_12290__bF_buf0) );
	BUFX4 BUFX4_742 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf5) );
	BUFX4 BUFX4_743 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf4) );
	BUFX4 BUFX4_744 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf3) );
	BUFX4 BUFX4_745 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf2) );
	BUFX4 BUFX4_746 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf1) );
	BUFX4 BUFX4_747 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .Y(_8417__bF_buf0) );
	BUFX4 BUFX4_748 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf8) );
	BUFX4 BUFX4_749 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf7) );
	BUFX4 BUFX4_750 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf6) );
	BUFX4 BUFX4_751 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf5) );
	BUFX4 BUFX4_752 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf4) );
	BUFX4 BUFX4_753 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf3) );
	BUFX4 BUFX4_754 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf2) );
	BUFX4 BUFX4_755 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf1) );
	BUFX4 BUFX4_756 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8616__bF_buf0) );
	BUFX4 BUFX4_757 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf42) );
	BUFX4 BUFX4_758 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf41) );
	BUFX4 BUFX4_759 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf40) );
	BUFX4 BUFX4_760 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf39) );
	BUFX4 BUFX4_761 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf38) );
	BUFX4 BUFX4_762 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf37) );
	BUFX4 BUFX4_763 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf36) );
	BUFX4 BUFX4_764 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf35) );
	BUFX4 BUFX4_765 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf34) );
	BUFX4 BUFX4_766 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf33) );
	BUFX4 BUFX4_767 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf32) );
	BUFX4 BUFX4_768 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf31) );
	BUFX4 BUFX4_769 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf30) );
	BUFX4 BUFX4_770 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf29) );
	BUFX4 BUFX4_771 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf28) );
	BUFX4 BUFX4_772 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf27) );
	BUFX4 BUFX4_773 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf26) );
	BUFX4 BUFX4_774 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf25) );
	BUFX4 BUFX4_775 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf24) );
	BUFX4 BUFX4_776 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf23) );
	BUFX4 BUFX4_777 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf22) );
	BUFX4 BUFX4_778 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf21) );
	BUFX4 BUFX4_779 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf20) );
	BUFX4 BUFX4_780 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf19) );
	BUFX4 BUFX4_781 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf18) );
	BUFX4 BUFX4_782 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf17) );
	BUFX4 BUFX4_783 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf16) );
	BUFX4 BUFX4_784 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf15) );
	BUFX4 BUFX4_785 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf14) );
	BUFX4 BUFX4_786 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf13) );
	BUFX4 BUFX4_787 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf12) );
	BUFX4 BUFX4_788 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf11) );
	BUFX4 BUFX4_789 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf10) );
	BUFX4 BUFX4_790 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf9) );
	BUFX4 BUFX4_791 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf8) );
	BUFX4 BUFX4_792 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf7) );
	BUFX4 BUFX4_793 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf6) );
	BUFX4 BUFX4_794 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf4), .Y(_6879__bF_buf5) );
	BUFX4 BUFX4_795 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf3), .Y(_6879__bF_buf4) );
	BUFX4 BUFX4_796 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf2), .Y(_6879__bF_buf3) );
	BUFX4 BUFX4_797 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf1), .Y(_6879__bF_buf2) );
	BUFX4 BUFX4_798 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf0), .Y(_6879__bF_buf1) );
	BUFX4 BUFX4_799 ( .gnd(gnd), .vdd(vdd), .A(_6879__hier0_bF_buf5), .Y(_6879__bF_buf0) );
	BUFX4 BUFX4_800 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf5) );
	BUFX4 BUFX4_801 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf4) );
	BUFX4 BUFX4_802 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf3) );
	BUFX4 BUFX4_803 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf2) );
	BUFX4 BUFX4_804 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf1) );
	BUFX4 BUFX4_805 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .Y(_8111__bF_buf0) );
	BUFX4 BUFX4_806 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_14789__bF_buf4) );
	BUFX4 BUFX4_807 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_14789__bF_buf3) );
	BUFX4 BUFX4_808 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_14789__bF_buf2) );
	BUFX4 BUFX4_809 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_14789__bF_buf1) );
	BUFX4 BUFX4_810 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_14789__bF_buf0) );
	BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_), .Y(biu_ins_29_bF_buf3) );
	BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_), .Y(biu_ins_29_bF_buf2) );
	BUFX4 BUFX4_811 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_), .Y(biu_ins_29_bF_buf1) );
	BUFX4 BUFX4_812 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_), .Y(biu_ins_29_bF_buf0) );
	BUFX4 BUFX4_813 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf7) );
	BUFX4 BUFX4_814 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf6) );
	BUFX4 BUFX4_815 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf5) );
	BUFX4 BUFX4_816 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf4) );
	BUFX4 BUFX4_817 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf3) );
	BUFX4 BUFX4_818 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf2) );
	BUFX4 BUFX4_819 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf1) );
	BUFX4 BUFX4_820 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11158__bF_buf0) );
	BUFX4 BUFX4_821 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .Y(_1379__bF_buf4) );
	BUFX4 BUFX4_822 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .Y(_1379__bF_buf3) );
	BUFX4 BUFX4_823 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .Y(_1379__bF_buf2) );
	BUFX4 BUFX4_824 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .Y(_1379__bF_buf1) );
	BUFX4 BUFX4_825 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .Y(_1379__bF_buf0) );
	BUFX4 BUFX4_826 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .Y(_14321__bF_buf3) );
	BUFX4 BUFX4_827 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .Y(_14321__bF_buf2) );
	BUFX4 BUFX4_828 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .Y(_14321__bF_buf1) );
	BUFX4 BUFX4_829 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .Y(_14321__bF_buf0) );
	BUFX4 BUFX4_830 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .Y(_9095__bF_buf4) );
	BUFX4 BUFX4_831 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .Y(_9095__bF_buf3) );
	BUFX4 BUFX4_832 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .Y(_9095__bF_buf2) );
	BUFX4 BUFX4_833 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .Y(_9095__bF_buf1) );
	BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .Y(_9095__bF_buf0) );
	BUFX4 BUFX4_834 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf15) );
	BUFX4 BUFX4_835 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf14) );
	BUFX4 BUFX4_836 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf13) );
	BUFX4 BUFX4_837 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf12) );
	BUFX4 BUFX4_838 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf11) );
	BUFX4 BUFX4_839 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf10) );
	BUFX4 BUFX4_840 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf9) );
	BUFX4 BUFX4_841 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf8) );
	BUFX4 BUFX4_842 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf7) );
	BUFX4 BUFX4_843 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf6) );
	BUFX4 BUFX4_844 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf5) );
	BUFX4 BUFX4_845 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf4) );
	BUFX4 BUFX4_846 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf3) );
	BUFX4 BUFX4_847 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf2) );
	BUFX4 BUFX4_848 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf1) );
	BUFX4 BUFX4_849 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3111__bF_buf0) );
	BUFX4 BUFX4_850 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_), .Y(addr_csr_21_bF_buf3) );
	BUFX4 BUFX4_851 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_), .Y(addr_csr_21_bF_buf2) );
	BUFX4 BUFX4_852 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_), .Y(addr_csr_21_bF_buf1) );
	BUFX4 BUFX4_853 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_), .Y(addr_csr_21_bF_buf0) );
	BUFX4 BUFX4_854 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf7) );
	BUFX4 BUFX4_855 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf6) );
	BUFX4 BUFX4_856 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf5) );
	BUFX4 BUFX4_857 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf4) );
	BUFX4 BUFX4_858 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf3) );
	BUFX4 BUFX4_859 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf2) );
	BUFX4 BUFX4_860 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf1) );
	BUFX4 BUFX4_861 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .Y(_4910__bF_buf0) );
	BUFX4 BUFX4_862 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .Y(_9234__bF_buf3) );
	BUFX4 BUFX4_863 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .Y(_9234__bF_buf2) );
	BUFX4 BUFX4_864 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .Y(_9234__bF_buf1) );
	BUFX4 BUFX4_865 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .Y(_9234__bF_buf0) );
	BUFX4 BUFX4_866 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .Y(_9162__bF_buf3) );
	BUFX4 BUFX4_867 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .Y(_9162__bF_buf2) );
	BUFX4 BUFX4_868 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .Y(_9162__bF_buf1) );
	BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .Y(_9162__bF_buf0) );
	BUFX4 BUFX4_869 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .Y(_2541__bF_buf4) );
	BUFX4 BUFX4_870 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .Y(_2541__bF_buf3) );
	BUFX4 BUFX4_871 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .Y(_2541__bF_buf2) );
	BUFX4 BUFX4_872 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .Y(_2541__bF_buf1) );
	BUFX4 BUFX4_873 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .Y(_2541__bF_buf0) );
	BUFX4 BUFX4_874 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(_2511__bF_buf4) );
	BUFX4 BUFX4_875 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(_2511__bF_buf3) );
	BUFX4 BUFX4_876 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(_2511__bF_buf2) );
	BUFX4 BUFX4_877 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(_2511__bF_buf1) );
	BUFX4 BUFX4_878 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(_2511__bF_buf0) );
	BUFX4 BUFX4_879 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf5) );
	BUFX4 BUFX4_880 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf4) );
	BUFX4 BUFX4_881 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf3) );
	BUFX4 BUFX4_882 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf2) );
	BUFX4 BUFX4_883 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf1) );
	BUFX4 BUFX4_884 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf0) );
	BUFX4 BUFX4_885 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_35__bF_buf3) );
	BUFX4 BUFX4_886 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_35__bF_buf2) );
	BUFX4 BUFX4_887 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_35__bF_buf1) );
	BUFX4 BUFX4_888 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_35__bF_buf0) );
	BUFX4 BUFX4_889 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf6) );
	BUFX4 BUFX4_890 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf5) );
	BUFX4 BUFX4_891 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf4) );
	BUFX4 BUFX4_892 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf3) );
	BUFX4 BUFX4_893 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf2) );
	BUFX4 BUFX4_894 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf1) );
	BUFX4 BUFX4_895 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .Y(_7594__bF_buf0) );
	BUFX4 BUFX4_896 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6193__bF_buf4) );
	BUFX4 BUFX4_897 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6193__bF_buf3) );
	BUFX4 BUFX4_898 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6193__bF_buf2) );
	BUFX4 BUFX4_899 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6193__bF_buf1) );
	BUFX4 BUFX4_900 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6193__bF_buf0) );
	BUFX4 BUFX4_901 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .Y(_7962__bF_buf4) );
	BUFX4 BUFX4_902 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .Y(_7962__bF_buf3) );
	BUFX4 BUFX4_903 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .Y(_7962__bF_buf2) );
	BUFX4 BUFX4_904 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .Y(_7962__bF_buf1) );
	BUFX4 BUFX4_905 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .Y(_7962__bF_buf0) );
	BUFX4 BUFX4_906 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .Y(_6392__bF_buf4) );
	BUFX4 BUFX4_907 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .Y(_6392__bF_buf3) );
	BUFX4 BUFX4_908 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .Y(_6392__bF_buf2) );
	BUFX4 BUFX4_909 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .Y(_6392__bF_buf1) );
	BUFX4 BUFX4_910 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .Y(_6392__bF_buf0) );
	BUFX4 BUFX4_911 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf10) );
	BUFX4 BUFX4_912 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf9) );
	BUFX4 BUFX4_913 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf8) );
	BUFX4 BUFX4_914 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf7) );
	BUFX4 BUFX4_915 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf6) );
	BUFX4 BUFX4_916 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf5) );
	BUFX4 BUFX4_917 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf4) );
	BUFX4 BUFX4_918 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf3) );
	BUFX4 BUFX4_919 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf2) );
	BUFX4 BUFX4_920 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf1) );
	BUFX4 BUFX4_921 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3109__bF_buf0) );
	BUFX4 BUFX4_922 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .Y(_13478__bF_buf4) );
	BUFX4 BUFX4_923 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .Y(_13478__bF_buf3) );
	BUFX4 BUFX4_924 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .Y(_13478__bF_buf2) );
	BUFX4 BUFX4_925 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .Y(_13478__bF_buf1) );
	BUFX4 BUFX4_926 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .Y(_13478__bF_buf0) );
	BUFX4 BUFX4_927 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf3) );
	BUFX4 BUFX4_928 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf2) );
	BUFX4 BUFX4_929 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf1) );
	BUFX4 BUFX4_930 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf0) );
	BUFX4 BUFX4_931 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_), .Y(addr_csr_19_bF_buf3) );
	BUFX4 BUFX4_932 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_), .Y(addr_csr_19_bF_buf2) );
	BUFX4 BUFX4_933 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_), .Y(addr_csr_19_bF_buf1) );
	BUFX4 BUFX4_934 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_), .Y(addr_csr_19_bF_buf0) );
	BUFX4 BUFX4_935 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6591__bF_buf4) );
	BUFX4 BUFX4_936 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6591__bF_buf3) );
	BUFX4 BUFX4_937 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6591__bF_buf2) );
	BUFX4 BUFX4_938 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6591__bF_buf1) );
	BUFX4 BUFX4_939 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6591__bF_buf0) );
	BUFX4 BUFX4_940 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf13) );
	BUFX4 BUFX4_941 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf12) );
	BUFX4 BUFX4_942 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf11) );
	BUFX4 BUFX4_943 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf10) );
	BUFX4 BUFX4_944 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf9) );
	BUFX4 BUFX4_945 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf8) );
	BUFX4 BUFX4_946 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf7) );
	BUFX4 BUFX4_947 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf6) );
	BUFX4 BUFX4_948 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf5) );
	BUFX4 BUFX4_949 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf4) );
	BUFX4 BUFX4_950 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf3) );
	BUFX4 BUFX4_951 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf2) );
	BUFX4 BUFX4_952 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf1) );
	BUFX4 BUFX4_953 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_4896__bF_buf0) );
	BUFX4 BUFX4_954 ( .gnd(gnd), .vdd(vdd), .A(_14916_), .Y(_14916__bF_buf3) );
	BUFX4 BUFX4_955 ( .gnd(gnd), .vdd(vdd), .A(_14916_), .Y(_14916__bF_buf2) );
	BUFX4 BUFX4_956 ( .gnd(gnd), .vdd(vdd), .A(_14916_), .Y(_14916__bF_buf1) );
	BUFX4 BUFX4_957 ( .gnd(gnd), .vdd(vdd), .A(_14916_), .Y(_14916__bF_buf0) );
	BUFX4 BUFX4_958 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .Y(_2539__bF_buf4) );
	BUFX4 BUFX4_959 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .Y(_2539__bF_buf3) );
	BUFX4 BUFX4_960 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .Y(_2539__bF_buf2) );
	BUFX4 BUFX4_961 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .Y(_2539__bF_buf1) );
	BUFX4 BUFX4_962 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .Y(_2539__bF_buf0) );
	BUFX4 BUFX4_963 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2509__bF_buf4) );
	BUFX4 BUFX4_964 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2509__bF_buf3) );
	BUFX4 BUFX4_965 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2509__bF_buf2) );
	BUFX4 BUFX4_966 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2509__bF_buf1) );
	BUFX4 BUFX4_967 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2509__bF_buf0) );
	BUFX4 BUFX4_968 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf4) );
	BUFX4 BUFX4_969 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf3) );
	BUFX4 BUFX4_970 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf2) );
	BUFX4 BUFX4_971 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf1) );
	BUFX4 BUFX4_972 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf0) );
	BUFX4 BUFX4_973 ( .gnd(gnd), .vdd(vdd), .A(_856_), .Y(_856__bF_buf3) );
	BUFX4 BUFX4_974 ( .gnd(gnd), .vdd(vdd), .A(_856_), .Y(_856__bF_buf2) );
	BUFX4 BUFX4_975 ( .gnd(gnd), .vdd(vdd), .A(_856_), .Y(_856__bF_buf1) );
	BUFX4 BUFX4_976 ( .gnd(gnd), .vdd(vdd), .A(_856_), .Y(_856__bF_buf0) );
	BUFX4 BUFX4_977 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_224__bF_buf4) );
	BUFX4 BUFX4_978 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_224__bF_buf3) );
	BUFX4 BUFX4_979 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_224__bF_buf2) );
	BUFX4 BUFX4_980 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_224__bF_buf1) );
	BUFX4 BUFX4_981 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_224__bF_buf0) );
	BUFX4 BUFX4_982 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf12) );
	BUFX4 BUFX4_983 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf11) );
	BUFX4 BUFX4_984 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf10) );
	BUFX4 BUFX4_985 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf9) );
	BUFX4 BUFX4_986 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf8) );
	BUFX4 BUFX4_987 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf7) );
	BUFX4 BUFX4_988 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf6) );
	BUFX4 BUFX4_989 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf5) );
	BUFX4 BUFX4_990 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf4) );
	BUFX4 BUFX4_991 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf3) );
	BUFX4 BUFX4_992 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf2) );
	BUFX4 BUFX4_993 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf1) );
	BUFX4 BUFX4_994 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .Y(_2696__bF_buf0) );
	BUFX4 BUFX4_995 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf9) );
	BUFX4 BUFX4_996 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf8) );
	BUFX4 BUFX4_997 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf7) );
	BUFX4 BUFX4_998 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf6) );
	BUFX4 BUFX4_999 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf5) );
	BUFX4 BUFX4_1000 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf4) );
	BUFX4 BUFX4_1001 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf3) );
	BUFX4 BUFX4_1002 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf2) );
	BUFX4 BUFX4_1003 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf1) );
	BUFX4 BUFX4_1004 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .Y(_4903__bF_buf0) );
	BUFX4 BUFX4_1005 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_), .Y(biu_exce_chk_statu_biu_6_bF_buf3) );
	BUFX4 BUFX4_1006 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_), .Y(biu_exce_chk_statu_biu_6_bF_buf2) );
	BUFX4 BUFX4_1007 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_), .Y(biu_exce_chk_statu_biu_6_bF_buf1) );
	BUFX4 BUFX4_1008 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_), .Y(biu_exce_chk_statu_biu_6_bF_buf0) );
	BUFX4 BUFX4_1009 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf7) );
	BUFX4 BUFX4_1010 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf6) );
	BUFX4 BUFX4_1011 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf5) );
	BUFX4 BUFX4_1012 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf4) );
	BUFX4 BUFX4_1013 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf3) );
	BUFX4 BUFX4_1014 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf2) );
	BUFX4 BUFX4_1015 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf1) );
	BUFX4 BUFX4_1016 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4891__bF_buf0) );
	BUFX4 BUFX4_1017 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .Y(_6059__bF_buf4) );
	BUFX4 BUFX4_1018 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .Y(_6059__bF_buf3) );
	BUFX4 BUFX4_1019 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .Y(_6059__bF_buf2) );
	BUFX4 BUFX4_1020 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .Y(_6059__bF_buf1) );
	BUFX4 BUFX4_1021 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .Y(_6059__bF_buf0) );
	BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp), .Y(csr_gpr_iu_ins_dec_subp_bF_buf3) );
	BUFX4 BUFX4_1022 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp), .Y(csr_gpr_iu_ins_dec_subp_bF_buf2) );
	BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp), .Y(csr_gpr_iu_ins_dec_subp_bF_buf1) );
	BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp), .Y(csr_gpr_iu_ins_dec_subp_bF_buf0) );
	BUFX4 BUFX4_1023 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_28__bF_buf3) );
	BUFX4 BUFX4_1024 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_28__bF_buf2) );
	BUFX4 BUFX4_1025 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_28__bF_buf1) );
	BUFX4 BUFX4_1026 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_28__bF_buf0) );
	BUFX4 BUFX4_1027 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .Y(_11412__bF_buf3) );
	BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .Y(_11412__bF_buf2) );
	BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .Y(_11412__bF_buf1) );
	BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .Y(_11412__bF_buf0) );
	BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf3) );
	BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf2) );
	BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf1) );
	BUFX4 BUFX4_1028 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf0) );
	BUFX4 BUFX4_1029 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_), .Y(biu_biu_data_out_7_bF_buf3) );
	BUFX4 BUFX4_1030 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_), .Y(biu_biu_data_out_7_bF_buf2) );
	BUFX4 BUFX4_1031 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_), .Y(biu_biu_data_out_7_bF_buf1) );
	BUFX4 BUFX4_1032 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_), .Y(biu_biu_data_out_7_bF_buf0) );
	BUFX4 BUFX4_1033 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_7323__bF_buf3) );
	BUFX4 BUFX4_1034 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_7323__bF_buf2) );
	BUFX4 BUFX4_1035 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_7323__bF_buf1) );
	BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_7323__bF_buf0) );
	BUFX4 BUFX4_1036 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf7) );
	BUFX4 BUFX4_1037 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf6) );
	BUFX4 BUFX4_1038 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf5) );
	BUFX4 BUFX4_1039 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf4) );
	BUFX4 BUFX4_1040 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf3) );
	BUFX4 BUFX4_1041 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf2) );
	BUFX4 BUFX4_1042 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf1) );
	BUFX4 BUFX4_1043 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal), .Y(csr_gpr_iu_ins_dec_jal_bF_buf0) );
	BUFX4 BUFX4_1044 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf5) );
	BUFX4 BUFX4_1045 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf4) );
	BUFX4 BUFX4_1046 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf3) );
	BUFX4 BUFX4_1047 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf2) );
	BUFX4 BUFX4_1048 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf1) );
	BUFX4 BUFX4_1049 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3127__bF_buf0) );
	BUFX4 BUFX4_1050 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf6) );
	BUFX4 BUFX4_1051 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf5) );
	BUFX4 BUFX4_1052 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf4) );
	BUFX4 BUFX4_1053 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf3) );
	BUFX4 BUFX4_1054 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf2) );
	BUFX4 BUFX4_1055 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf1) );
	BUFX4 BUFX4_1056 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13466__bF_buf0) );
	BUFX4 BUFX4_1057 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf5) );
	BUFX4 BUFX4_1058 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf4) );
	BUFX4 BUFX4_1059 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf3) );
	BUFX4 BUFX4_1060 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf2) );
	BUFX4 BUFX4_1061 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf1) );
	BUFX4 BUFX4_1062 ( .gnd(gnd), .vdd(vdd), .A(_13695_), .Y(_13695__bF_buf0) );
	BUFX4 BUFX4_1063 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .Y(_6820__bF_buf3) );
	BUFX4 BUFX4_1064 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .Y(_6820__bF_buf2) );
	BUFX4 BUFX4_1065 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .Y(_6820__bF_buf1) );
	BUFX4 BUFX4_1066 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .Y(_6820__bF_buf0) );
	BUFX4 BUFX4_1067 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .Y(_2527__bF_buf4) );
	BUFX4 BUFX4_1068 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .Y(_2527__bF_buf3) );
	BUFX4 BUFX4_1069 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .Y(_2527__bF_buf2) );
	BUFX4 BUFX4_1070 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .Y(_2527__bF_buf1) );
	BUFX4 BUFX4_1071 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .Y(_2527__bF_buf0) );
	BUFX4 BUFX4_1072 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf6) );
	BUFX4 BUFX4_1073 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf5) );
	BUFX4 BUFX4_1074 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf4) );
	BUFX4 BUFX4_1075 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf3) );
	BUFX4 BUFX4_1076 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf2) );
	BUFX4 BUFX4_1077 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf1) );
	BUFX4 BUFX4_1078 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_645__bF_buf0) );
	BUFX4 BUFX4_1079 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf5) );
	BUFX4 BUFX4_1080 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf4) );
	BUFX4 BUFX4_1081 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf3) );
	BUFX4 BUFX4_1082 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf2) );
	BUFX4 BUFX4_1083 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf1) );
	BUFX4 BUFX4_1084 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .Y(_1228__bF_buf0) );
	BUFX4 BUFX4_1085 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb), .Y(biu_ahb_statu_ahb_bF_buf4) );
	BUFX4 BUFX4_1086 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb), .Y(biu_ahb_statu_ahb_bF_buf3) );
	BUFX4 BUFX4_1087 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb), .Y(biu_ahb_statu_ahb_bF_buf2) );
	BUFX4 BUFX4_1088 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb), .Y(biu_ahb_statu_ahb_bF_buf1) );
	BUFX4 BUFX4_1089 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb), .Y(biu_ahb_statu_ahb_bF_buf0) );
	BUFX4 BUFX4_1090 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_), .Y(biu_ins_30_bF_buf3) );
	BUFX4 BUFX4_1091 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_), .Y(biu_ins_30_bF_buf2) );
	BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_), .Y(biu_ins_30_bF_buf1) );
	BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_), .Y(biu_ins_30_bF_buf0) );
	BUFX4 BUFX4_1092 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .Y(_12132__bF_buf3) );
	BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .Y(_12132__bF_buf2) );
	BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .Y(_12132__bF_buf1) );
	BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .Y(_12132__bF_buf0) );
	BUFX4 BUFX4_1093 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .Y(_2624__bF_buf4) );
	BUFX4 BUFX4_1094 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .Y(_2624__bF_buf3) );
	BUFX4 BUFX4_1095 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .Y(_2624__bF_buf2) );
	BUFX4 BUFX4_1096 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .Y(_2624__bF_buf1) );
	BUFX4 BUFX4_1097 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .Y(_2624__bF_buf0) );
	BUFX4 BUFX4_1098 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf4) );
	BUFX4 BUFX4_1099 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf3) );
	BUFX4 BUFX4_1100 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf2) );
	BUFX4 BUFX4_1101 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf1) );
	BUFX4 BUFX4_1102 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf0) );
	BUFX4 BUFX4_1103 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .Y(_13459__bF_buf4) );
	BUFX4 BUFX4_1104 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .Y(_13459__bF_buf3) );
	BUFX4 BUFX4_1105 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .Y(_13459__bF_buf2) );
	BUFX4 BUFX4_1106 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .Y(_13459__bF_buf1) );
	BUFX4 BUFX4_1107 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .Y(_13459__bF_buf0) );
	BUFX4 BUFX4_1108 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_2__bF_buf3) );
	BUFX4 BUFX4_1109 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_2__bF_buf2) );
	BUFX4 BUFX4_1110 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_2__bF_buf1) );
	BUFX4 BUFX4_1111 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_2__bF_buf0) );
	BUFX4 BUFX4_1112 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_), .Y(biu_ins_28_bF_buf3) );
	BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_), .Y(biu_ins_28_bF_buf2) );
	BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_), .Y(biu_ins_28_bF_buf1) );
	BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_), .Y(biu_ins_28_bF_buf0) );
	BUFX4 BUFX4_1113 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_14825__bF_buf4) );
	BUFX4 BUFX4_1114 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_14825__bF_buf3) );
	BUFX4 BUFX4_1115 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_14825__bF_buf2) );
	BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_14825__bF_buf1) );
	BUFX4 BUFX4_1116 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_14825__bF_buf0) );
	BUFX4 BUFX4_1117 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_837__bF_buf3) );
	BUFX4 BUFX4_1118 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_837__bF_buf2) );
	BUFX4 BUFX4_1119 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_837__bF_buf1) );
	BUFX4 BUFX4_1120 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_837__bF_buf0) );
	BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .Y(_13454__bF_buf4) );
	BUFX4 BUFX4_1121 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .Y(_13454__bF_buf3) );
	BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .Y(_13454__bF_buf2) );
	BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .Y(_13454__bF_buf1) );
	BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .Y(_13454__bF_buf0) );
	BUFX4 BUFX4_1122 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_), .Y(addr_csr_25_bF_buf3) );
	BUFX4 BUFX4_1123 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_), .Y(addr_csr_25_bF_buf2) );
	BUFX4 BUFX4_1124 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_), .Y(addr_csr_25_bF_buf1) );
	BUFX4 BUFX4_1125 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_), .Y(addr_csr_25_bF_buf0) );
	BUFX4 BUFX4_1126 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .Y(_11127__bF_buf4) );
	BUFX4 BUFX4_1127 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .Y(_11127__bF_buf3) );
	BUFX4 BUFX4_1128 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .Y(_11127__bF_buf2) );
	BUFX4 BUFX4_1129 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .Y(_11127__bF_buf1) );
	BUFX4 BUFX4_1130 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .Y(_11127__bF_buf0) );
	BUFX4 BUFX4_1131 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf6) );
	BUFX4 BUFX4_1132 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf5) );
	BUFX4 BUFX4_1133 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf4) );
	BUFX4 BUFX4_1134 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf3) );
	BUFX4 BUFX4_1135 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf2) );
	BUFX4 BUFX4_1136 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf1) );
	BUFX4 BUFX4_1137 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .Y(_9268__bF_buf0) );
	BUFX4 BUFX4_1138 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2545__bF_buf4) );
	BUFX4 BUFX4_1139 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2545__bF_buf3) );
	BUFX4 BUFX4_1140 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2545__bF_buf2) );
	BUFX4 BUFX4_1141 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2545__bF_buf1) );
	BUFX4 BUFX4_1142 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2545__bF_buf0) );
	BUFX4 BUFX4_1143 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .Y(_2515__bF_buf4) );
	BUFX4 BUFX4_1144 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .Y(_2515__bF_buf3) );
	BUFX4 BUFX4_1145 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .Y(_2515__bF_buf2) );
	BUFX4 BUFX4_1146 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .Y(_2515__bF_buf1) );
	BUFX4 BUFX4_1147 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .Y(_2515__bF_buf0) );
	BUFX4 BUFX4_1148 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf5) );
	BUFX4 BUFX4_1149 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf4) );
	BUFX4 BUFX4_1150 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf3) );
	BUFX4 BUFX4_1151 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf2) );
	BUFX4 BUFX4_1152 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf1) );
	BUFX4 BUFX4_1153 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .Y(_9094__bF_buf0) );
	BUFX4 BUFX4_1154 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf7) );
	BUFX4 BUFX4_1155 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf6) );
	BUFX4 BUFX4_1156 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf5) );
	BUFX4 BUFX4_1157 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf4) );
	BUFX4 BUFX4_1158 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf3) );
	BUFX4 BUFX4_1159 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf2) );
	BUFX4 BUFX4_1160 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf1) );
	BUFX4 BUFX4_1161 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2473__bF_buf0) );
	BUFX4 BUFX4_1162 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf13) );
	BUFX4 BUFX4_1163 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf12) );
	BUFX4 BUFX4_1164 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf11) );
	BUFX4 BUFX4_1165 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf10) );
	BUFX4 BUFX4_1166 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf9) );
	BUFX4 BUFX4_1167 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf8) );
	BUFX4 BUFX4_1168 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf7) );
	BUFX4 BUFX4_1169 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf6) );
	BUFX4 BUFX4_1170 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf5) );
	BUFX4 BUFX4_1171 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf4) );
	BUFX4 BUFX4_1172 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf3) );
	BUFX4 BUFX4_1173 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf2) );
	BUFX4 BUFX4_1174 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf1) );
	BUFX4 BUFX4_1175 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .Y(_3110__bF_buf0) );
	BUFX4 BUFX4_1176 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_), .Y(biu_mmu_pte_new_7_bF_buf4) );
	BUFX4 BUFX4_1177 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_), .Y(biu_mmu_pte_new_7_bF_buf3) );
	BUFX4 BUFX4_1178 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_), .Y(biu_mmu_pte_new_7_bF_buf2) );
	BUFX4 BUFX4_1179 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_), .Y(biu_mmu_pte_new_7_bF_buf1) );
	BUFX4 BUFX4_1180 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_), .Y(biu_mmu_pte_new_7_bF_buf0) );
	BUFX4 BUFX4_1181 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .Y(_7309__bF_buf3) );
	BUFX4 BUFX4_1182 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .Y(_7309__bF_buf2) );
	BUFX4 BUFX4_1183 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .Y(_7309__bF_buf1) );
	BUFX4 BUFX4_1184 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .Y(_7309__bF_buf0) );
	BUFX4 BUFX4_1185 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf5) );
	BUFX4 BUFX4_1186 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf4) );
	BUFX4 BUFX4_1187 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf3) );
	BUFX4 BUFX4_1188 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf2) );
	BUFX4 BUFX4_1189 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf1) );
	BUFX4 BUFX4_1190 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .Y(_8235__bF_buf0) );
	BUFX4 BUFX4_1191 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9161__bF_buf4) );
	BUFX4 BUFX4_1192 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9161__bF_buf3) );
	BUFX4 BUFX4_1193 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9161__bF_buf2) );
	BUFX4 BUFX4_1194 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9161__bF_buf1) );
	BUFX4 BUFX4_1195 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9161__bF_buf0) );
	BUFX4 BUFX4_1196 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf14) );
	BUFX4 BUFX4_1197 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf13) );
	BUFX4 BUFX4_1198 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf12) );
	BUFX4 BUFX4_1199 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf11) );
	BUFX4 BUFX4_1200 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf10) );
	BUFX4 BUFX4_1201 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf9) );
	BUFX4 BUFX4_1202 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf8) );
	BUFX4 BUFX4_1203 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf7) );
	BUFX4 BUFX4_1204 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf6) );
	BUFX4 BUFX4_1205 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf5) );
	BUFX4 BUFX4_1206 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf4) );
	BUFX4 BUFX4_1207 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf3) );
	BUFX4 BUFX4_1208 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf2) );
	BUFX4 BUFX4_1209 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf1) );
	BUFX4 BUFX4_1210 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .Y(_7304__bF_buf0) );
	BUFX4 BUFX4_1211 ( .gnd(gnd), .vdd(vdd), .A(amoxor), .Y(amoxor_bF_buf3) );
	BUFX4 BUFX4_1212 ( .gnd(gnd), .vdd(vdd), .A(amoxor), .Y(amoxor_bF_buf2) );
	BUFX4 BUFX4_1213 ( .gnd(gnd), .vdd(vdd), .A(amoxor), .Y(amoxor_bF_buf1) );
	BUFX4 BUFX4_1214 ( .gnd(gnd), .vdd(vdd), .A(amoxor), .Y(amoxor_bF_buf0) );
	BUFX4 BUFX4_1215 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf10) );
	BUFX4 BUFX4_1216 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf9) );
	BUFX4 BUFX4_1217 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf8) );
	BUFX4 BUFX4_1218 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf7) );
	BUFX4 BUFX4_1219 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf6) );
	BUFX4 BUFX4_1220 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf5) );
	BUFX4 BUFX4_1221 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf4) );
	BUFX4 BUFX4_1222 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf3) );
	BUFX4 BUFX4_1223 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf2) );
	BUFX4 BUFX4_1224 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf1) );
	BUFX4 BUFX4_1225 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_4895__bF_buf0) );
	BUFX4 BUFX4_1226 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .Y(_2797__bF_buf4) );
	BUFX4 BUFX4_1227 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .Y(_2797__bF_buf3) );
	BUFX4 BUFX4_1228 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .Y(_2797__bF_buf2) );
	BUFX4 BUFX4_1229 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .Y(_2797__bF_buf1) );
	BUFX4 BUFX4_1230 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .Y(_2797__bF_buf0) );
	BUFX4 BUFX4_1231 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf7) );
	BUFX4 BUFX4_1232 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf6) );
	BUFX4 BUFX4_1233 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf5) );
	BUFX4 BUFX4_1234 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf4) );
	BUFX4 BUFX4_1235 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf3) );
	BUFX4 BUFX4_1236 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf2) );
	BUFX4 BUFX4_1237 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf1) );
	BUFX4 BUFX4_1238 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_223__bF_buf0) );
	BUFX4 BUFX4_1239 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .Y(_13412__bF_buf4) );
	BUFX4 BUFX4_1240 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .Y(_13412__bF_buf3) );
	BUFX4 BUFX4_1241 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .Y(_13412__bF_buf2) );
	BUFX4 BUFX4_1242 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .Y(_13412__bF_buf1) );
	BUFX4 BUFX4_1243 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .Y(_13412__bF_buf0) );
	BUFX4 BUFX4_1244 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .Y(_2695__bF_buf4) );
	BUFX4 BUFX4_1245 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .Y(_2695__bF_buf3) );
	BUFX4 BUFX4_1246 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .Y(_2695__bF_buf2) );
	BUFX4 BUFX4_1247 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .Y(_2695__bF_buf1) );
	BUFX4 BUFX4_1248 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .Y(_2695__bF_buf0) );
	BUFX4 BUFX4_1249 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_), .Y(addr_csr_13_bF_buf3) );
	BUFX4 BUFX4_1250 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_), .Y(addr_csr_13_bF_buf2) );
	BUFX4 BUFX4_1251 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_), .Y(addr_csr_13_bF_buf1) );
	BUFX4 BUFX4_1252 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_), .Y(addr_csr_13_bF_buf0) );
	BUFX4 BUFX4_1253 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .Y(_2533__bF_buf4) );
	BUFX4 BUFX4_1254 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .Y(_2533__bF_buf3) );
	BUFX4 BUFX4_1255 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .Y(_2533__bF_buf2) );
	BUFX4 BUFX4_1256 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .Y(_2533__bF_buf1) );
	BUFX4 BUFX4_1257 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .Y(_2533__bF_buf0) );
	BUFX4 BUFX4_1258 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_2503__bF_buf4) );
	BUFX4 BUFX4_1259 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_2503__bF_buf3) );
	BUFX4 BUFX4_1260 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_2503__bF_buf2) );
	BUFX4 BUFX4_1261 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_2503__bF_buf1) );
	BUFX4 BUFX4_1262 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_2503__bF_buf0) );
	BUFX4 BUFX4_1263 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .Y(_2491__bF_buf4) );
	BUFX4 BUFX4_1264 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .Y(_2491__bF_buf3) );
	BUFX4 BUFX4_1265 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .Y(_2491__bF_buf2) );
	BUFX4 BUFX4_1266 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .Y(_2491__bF_buf1) );
	BUFX4 BUFX4_1267 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .Y(_2491__bF_buf0) );
	BUFX4 BUFX4_1268 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf8) );
	BUFX4 BUFX4_1269 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf7) );
	BUFX4 BUFX4_1270 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf6) );
	BUFX4 BUFX4_1271 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf5) );
	BUFX4 BUFX4_1272 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf4) );
	BUFX4 BUFX4_1273 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf3) );
	BUFX4 BUFX4_1274 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf2) );
	BUFX4 BUFX4_1275 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf1) );
	BUFX4 BUFX4_1276 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_2732__bF_buf0) );
	BUFX4 BUFX4_1277 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6359__bF_buf4) );
	BUFX4 BUFX4_1278 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6359__bF_buf3) );
	BUFX4 BUFX4_1279 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6359__bF_buf2) );
	BUFX4 BUFX4_1280 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6359__bF_buf1) );
	BUFX4 BUFX4_1281 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6359__bF_buf0) );
	BUFX4 BUFX4_1282 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_27__bF_buf3) );
	BUFX4 BUFX4_1283 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_27__bF_buf2) );
	BUFX4 BUFX4_1284 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_27__bF_buf1) );
	BUFX4 BUFX4_1285 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_27__bF_buf0) );
	BUFX4 BUFX4_1286 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9281__bF_buf3) );
	BUFX4 BUFX4_1287 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9281__bF_buf2) );
	BUFX4 BUFX4_1288 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9281__bF_buf1) );
	BUFX4 BUFX4_1289 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9281__bF_buf0) );
	BUFX4 BUFX4_1290 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf6) );
	BUFX4 BUFX4_1291 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf5) );
	BUFX4 BUFX4_1292 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf4) );
	BUFX4 BUFX4_1293 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf3) );
	BUFX4 BUFX4_1294 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf2) );
	BUFX4 BUFX4_1295 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf1) );
	BUFX4 BUFX4_1296 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .Y(_9251__bF_buf0) );
	BUFX4 BUFX4_1297 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf70) );
	BUFX4 BUFX4_1298 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf69) );
	BUFX4 BUFX4_1299 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf68) );
	BUFX4 BUFX4_1300 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf67) );
	BUFX4 BUFX4_1301 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf66) );
	BUFX4 BUFX4_1302 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf65) );
	BUFX4 BUFX4_1303 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf64) );
	BUFX4 BUFX4_1304 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf63) );
	BUFX4 BUFX4_1305 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf62) );
	BUFX4 BUFX4_1306 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf61) );
	BUFX4 BUFX4_1307 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf60) );
	BUFX4 BUFX4_1308 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf59) );
	BUFX4 BUFX4_1309 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf58) );
	BUFX4 BUFX4_1310 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf57) );
	BUFX4 BUFX4_1311 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf56) );
	BUFX4 BUFX4_1312 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf55) );
	BUFX4 BUFX4_1313 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf54) );
	BUFX4 BUFX4_1314 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf53) );
	BUFX4 BUFX4_1315 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf52) );
	BUFX4 BUFX4_1316 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf51) );
	BUFX4 BUFX4_1317 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf50) );
	BUFX4 BUFX4_1318 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf49) );
	BUFX4 BUFX4_1319 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf48) );
	BUFX4 BUFX4_1320 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf47) );
	BUFX4 BUFX4_1321 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf46) );
	BUFX4 BUFX4_1322 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf45) );
	BUFX4 BUFX4_1323 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf44) );
	BUFX4 BUFX4_1324 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf43) );
	BUFX4 BUFX4_1325 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf42) );
	BUFX4 BUFX4_1326 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf41) );
	BUFX4 BUFX4_1327 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf40) );
	BUFX4 BUFX4_1328 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf39) );
	BUFX4 BUFX4_1329 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf38) );
	BUFX4 BUFX4_1330 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf37) );
	BUFX4 BUFX4_1331 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf36) );
	BUFX4 BUFX4_1332 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf35) );
	BUFX4 BUFX4_1333 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf34) );
	BUFX4 BUFX4_1334 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf33) );
	BUFX4 BUFX4_1335 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf32) );
	BUFX4 BUFX4_1336 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf31) );
	BUFX4 BUFX4_1337 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf30) );
	BUFX4 BUFX4_1338 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf29) );
	BUFX4 BUFX4_1339 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf28) );
	BUFX4 BUFX4_1340 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf27) );
	BUFX4 BUFX4_1341 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf26) );
	BUFX4 BUFX4_1342 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf25) );
	BUFX4 BUFX4_1343 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf24) );
	BUFX4 BUFX4_1344 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf23) );
	BUFX4 BUFX4_1345 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf22) );
	BUFX4 BUFX4_1346 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf21) );
	BUFX4 BUFX4_1347 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf20) );
	BUFX4 BUFX4_1348 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf19) );
	BUFX4 BUFX4_1349 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf18) );
	BUFX4 BUFX4_1350 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf17) );
	BUFX4 BUFX4_1351 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf16) );
	BUFX4 BUFX4_1352 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf15) );
	BUFX4 BUFX4_1353 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf14) );
	BUFX4 BUFX4_1354 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf13) );
	BUFX4 BUFX4_1355 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf12) );
	BUFX4 BUFX4_1356 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf11) );
	BUFX4 BUFX4_1357 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf10) );
	BUFX4 BUFX4_1358 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf9) );
	BUFX4 BUFX4_1359 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf8) );
	BUFX4 BUFX4_1360 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf0), .Y(rst_bF_buf7) );
	BUFX4 BUFX4_1361 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf7), .Y(rst_bF_buf6) );
	BUFX4 BUFX4_1362 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf6), .Y(rst_bF_buf5) );
	BUFX4 BUFX4_1363 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf5), .Y(rst_bF_buf4) );
	BUFX4 BUFX4_1364 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf4), .Y(rst_bF_buf3) );
	BUFX4 BUFX4_1365 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf3), .Y(rst_bF_buf2) );
	BUFX4 BUFX4_1366 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf2), .Y(rst_bF_buf1) );
	BUFX4 BUFX4_1367 ( .gnd(gnd), .vdd(vdd), .A(rst_hier0_bF_buf1), .Y(rst_bF_buf0) );
	BUFX4 BUFX4_1368 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf5) );
	BUFX4 BUFX4_1369 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf4) );
	BUFX4 BUFX4_1370 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf3) );
	BUFX4 BUFX4_1371 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf2) );
	BUFX4 BUFX4_1372 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf1) );
	BUFX4 BUFX4_1373 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .Y(_7586__bF_buf0) );
	BUFX4 BUFX4_1374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf6) );
	BUFX4 BUFX4_1375 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf5) );
	BUFX4 BUFX4_1376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf4) );
	BUFX4 BUFX4_1377 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf3) );
	BUFX4 BUFX4_1378 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf2) );
	BUFX4 BUFX4_1379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf1) );
	BUFX4 BUFX4_1380 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_), .Y(csr_gpr_iu_cause_31_bF_buf0) );
	BUFX4 BUFX4_1381 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6558__bF_buf4) );
	BUFX4 BUFX4_1382 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6558__bF_buf3) );
	BUFX4 BUFX4_1383 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6558__bF_buf2) );
	BUFX4 BUFX4_1384 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6558__bF_buf1) );
	BUFX4 BUFX4_1385 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6558__bF_buf0) );
	BUFX4 BUFX4_1386 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .Y(_7424__bF_buf3) );
	BUFX4 BUFX4_1387 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .Y(_7424__bF_buf2) );
	BUFX4 BUFX4_1388 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .Y(_7424__bF_buf1) );
	BUFX4 BUFX4_1389 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .Y(_7424__bF_buf0) );
	BUFX4 BUFX4_1390 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf10) );
	BUFX4 BUFX4_1391 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf9) );
	BUFX4 BUFX4_1392 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf8) );
	BUFX4 BUFX4_1393 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf7) );
	BUFX4 BUFX4_1394 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf6) );
	BUFX4 BUFX4_1395 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf5) );
	BUFX4 BUFX4_1396 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf4) );
	BUFX4 BUFX4_1397 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf3) );
	BUFX4 BUFX4_1398 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf2) );
	BUFX4 BUFX4_1399 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf1) );
	BUFX4 BUFX4_1400 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_6426__bF_buf0) );
	BUFX4 BUFX4_1401 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .Y(_6125__bF_buf4) );
	BUFX4 BUFX4_1402 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .Y(_6125__bF_buf3) );
	BUFX4 BUFX4_1403 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .Y(_6125__bF_buf2) );
	BUFX4 BUFX4_1404 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .Y(_6125__bF_buf1) );
	BUFX4 BUFX4_1405 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .Y(_6125__bF_buf0) );
	BUFX4 BUFX4_1406 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(_8621__bF_buf4) );
	BUFX4 BUFX4_1407 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(_8621__bF_buf3) );
	BUFX4 BUFX4_1408 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(_8621__bF_buf2) );
	BUFX4 BUFX4_1409 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(_8621__bF_buf1) );
	BUFX4 BUFX4_1410 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(_8621__bF_buf0) );
	BUFX4 BUFX4_1411 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_7021__bF_buf4) );
	BUFX4 BUFX4_1412 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_7021__bF_buf3) );
	BUFX4 BUFX4_1413 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_7021__bF_buf2) );
	BUFX4 BUFX4_1414 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_7021__bF_buf1) );
	BUFX4 BUFX4_1415 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_7021__bF_buf0) );
	BUFX4 BUFX4_1416 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .Y(_3059__bF_buf4) );
	BUFX4 BUFX4_1417 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .Y(_3059__bF_buf3) );
	BUFX4 BUFX4_1418 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .Y(_3059__bF_buf2) );
	BUFX4 BUFX4_1419 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .Y(_3059__bF_buf1) );
	BUFX4 BUFX4_1420 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .Y(_3059__bF_buf0) );
	BUFX4 BUFX4_1421 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf6) );
	BUFX4 BUFX4_1422 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf5) );
	BUFX4 BUFX4_1423 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf4) );
	BUFX4 BUFX4_1424 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf3) );
	BUFX4 BUFX4_1425 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf2) );
	BUFX4 BUFX4_1426 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf1) );
	BUFX4 BUFX4_1427 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .Y(_13398__bF_buf0) );
	BUFX4 BUFX4_1428 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .Y(_14896__bF_buf4) );
	BUFX4 BUFX4_1429 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .Y(_14896__bF_buf3) );
	BUFX4 BUFX4_1430 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .Y(_14896__bF_buf2) );
	BUFX4 BUFX4_1431 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .Y(_14896__bF_buf1) );
	BUFX4 BUFX4_1432 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .Y(_14896__bF_buf0) );
	BUFX4 BUFX4_1433 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3156__bF_buf4) );
	BUFX4 BUFX4_1434 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3156__bF_buf3) );
	BUFX4 BUFX4_1435 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3156__bF_buf2) );
	BUFX4 BUFX4_1436 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3156__bF_buf1) );
	BUFX4 BUFX4_1437 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3156__bF_buf0) );
	BUFX4 BUFX4_1438 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .Y(_2489__bF_buf4) );
	BUFX4 BUFX4_1439 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .Y(_2489__bF_buf3) );
	BUFX4 BUFX4_1440 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .Y(_2489__bF_buf2) );
	BUFX4 BUFX4_1441 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .Y(_2489__bF_buf1) );
	BUFX4 BUFX4_1442 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .Y(_2489__bF_buf0) );
	BUFX4 BUFX4_1443 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf7) );
	BUFX4 BUFX4_1444 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf6) );
	BUFX4 BUFX4_1445 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf5) );
	BUFX4 BUFX4_1446 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf4) );
	BUFX4 BUFX4_1447 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf3) );
	BUFX4 BUFX4_1448 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf2) );
	BUFX4 BUFX4_1449 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf1) );
	BUFX4 BUFX4_1450 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .Y(_3126__bF_buf0) );
	BUFX4 BUFX4_1451 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf4) );
	BUFX4 BUFX4_1452 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf3) );
	BUFX4 BUFX4_1453 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf2) );
	BUFX4 BUFX4_1454 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf1) );
	BUFX4 BUFX4_1455 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf0) );
	BUFX4 BUFX4_1456 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2658__bF_buf4) );
	BUFX4 BUFX4_1457 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2658__bF_buf3) );
	BUFX4 BUFX4_1458 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2658__bF_buf2) );
	BUFX4 BUFX4_1459 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2658__bF_buf1) );
	BUFX4 BUFX4_1460 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2658__bF_buf0) );
	BUFX4 BUFX4_1461 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .Y(_13694__bF_buf4) );
	BUFX4 BUFX4_1462 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .Y(_13694__bF_buf3) );
	BUFX4 BUFX4_1463 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .Y(_13694__bF_buf2) );
	BUFX4 BUFX4_1464 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .Y(_13694__bF_buf1) );
	BUFX4 BUFX4_1465 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .Y(_13694__bF_buf0) );
	BUFX4 BUFX4_1466 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .Y(_14331__bF_buf3) );
	BUFX4 BUFX4_1467 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .Y(_14331__bF_buf2) );
	BUFX4 BUFX4_1468 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .Y(_14331__bF_buf1) );
	BUFX4 BUFX4_1469 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .Y(_14331__bF_buf0) );
	BUFX4 BUFX4_1470 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf5) );
	BUFX4 BUFX4_1471 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf4) );
	BUFX4 BUFX4_1472 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf3) );
	BUFX4 BUFX4_1473 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf2) );
	BUFX4 BUFX4_1474 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf1) );
	BUFX4 BUFX4_1475 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf0) );
	BUFX4 BUFX4_1476 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .Y(_12305__bF_buf4) );
	BUFX4 BUFX4_1477 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .Y(_12305__bF_buf3) );
	BUFX4 BUFX4_1478 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .Y(_12305__bF_buf2) );
	BUFX4 BUFX4_1479 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .Y(_12305__bF_buf1) );
	BUFX4 BUFX4_1480 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .Y(_12305__bF_buf0) );
	BUFX4 BUFX4_1481 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf12) );
	BUFX4 BUFX4_1482 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf11) );
	BUFX4 BUFX4_1483 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf10) );
	BUFX4 BUFX4_1484 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf9) );
	BUFX4 BUFX4_1485 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf8) );
	BUFX4 BUFX4_1486 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf7) );
	BUFX4 BUFX4_1487 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf6) );
	BUFX4 BUFX4_1488 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf5) );
	BUFX4 BUFX4_1489 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf4) );
	BUFX4 BUFX4_1490 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf3) );
	BUFX4 BUFX4_1491 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf2) );
	BUFX4 BUFX4_1492 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf1) );
	BUFX4 BUFX4_1493 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .Y(_2484__bF_buf0) );
	BUFX4 BUFX4_1494 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_), .Y(addr_csr_31_bF_buf3) );
	BUFX4 BUFX4_1495 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_), .Y(addr_csr_31_bF_buf2) );
	BUFX4 BUFX4_1496 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_), .Y(addr_csr_31_bF_buf1) );
	BUFX4 BUFX4_1497 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_), .Y(addr_csr_31_bF_buf0) );
	BUFX4 BUFX4_1498 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .Y(_2521__bF_buf4) );
	BUFX4 BUFX4_1499 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .Y(_2521__bF_buf3) );
	BUFX4 BUFX4_1500 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .Y(_2521__bF_buf2) );
	BUFX4 BUFX4_1501 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .Y(_2521__bF_buf1) );
	BUFX4 BUFX4_1502 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .Y(_2521__bF_buf0) );
	BUFX4 BUFX4_1503 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf5) );
	BUFX4 BUFX4_1504 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf4) );
	BUFX4 BUFX4_1505 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf3) );
	BUFX4 BUFX4_1506 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf2) );
	BUFX4 BUFX4_1507 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf1) );
	BUFX4 BUFX4_1508 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .Y(_1222__bF_buf0) );
	BUFX4 BUFX4_1509 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf5) );
	BUFX4 BUFX4_1510 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf4) );
	BUFX4 BUFX4_1511 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf3) );
	BUFX4 BUFX4_1512 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf2) );
	BUFX4 BUFX4_1513 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf1) );
	BUFX4 BUFX4_1514 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .Y(_8373__bF_buf0) );
	BUFX4 BUFX4_1515 ( .gnd(gnd), .vdd(vdd), .A(_13488_), .Y(_13488__bF_buf3) );
	BUFX4 BUFX4_1516 ( .gnd(gnd), .vdd(vdd), .A(_13488_), .Y(_13488__bF_buf2) );
	BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(_13488_), .Y(_13488__bF_buf1) );
	BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(_13488_), .Y(_13488__bF_buf0) );
	BUFX4 BUFX4_1517 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf8) );
	BUFX4 BUFX4_1518 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf7) );
	BUFX4 BUFX4_1519 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf6) );
	BUFX4 BUFX4_1520 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf5) );
	BUFX4 BUFX4_1521 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf4) );
	BUFX4 BUFX4_1522 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf3) );
	BUFX4 BUFX4_1523 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf2) );
	BUFX4 BUFX4_1524 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf1) );
	BUFX4 BUFX4_1525 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13458__bF_buf0) );
	BUFX4 BUFX4_1526 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_), .Y(biu_ins_27_bF_buf3) );
	BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_), .Y(biu_ins_27_bF_buf2) );
	BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_), .Y(biu_ins_27_bF_buf1) );
	BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_), .Y(biu_ins_27_bF_buf0) );
	BUFX4 BUFX4_1527 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_), .Y(addr_csr_29_bF_buf3) );
	BUFX4 BUFX4_1528 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_), .Y(addr_csr_29_bF_buf2) );
	BUFX4 BUFX4_1529 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_), .Y(addr_csr_29_bF_buf1) );
	BUFX4 BUFX4_1530 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_), .Y(addr_csr_29_bF_buf0) );
	BUFX4 BUFX4_1531 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf7) );
	BUFX4 BUFX4_1532 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf6) );
	BUFX4 BUFX4_1533 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf5) );
	BUFX4 BUFX4_1534 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf4) );
	BUFX4 BUFX4_1535 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf3) );
	BUFX4 BUFX4_1536 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf2) );
	BUFX4 BUFX4_1537 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf1) );
	BUFX4 BUFX4_1538 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .Y(_13687__bF_buf0) );
	BUFX4 BUFX4_1539 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf8) );
	BUFX4 BUFX4_1540 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf7) );
	BUFX4 BUFX4_1541 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf6) );
	BUFX4 BUFX4_1542 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf5) );
	BUFX4 BUFX4_1543 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf4) );
	BUFX4 BUFX4_1544 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf3) );
	BUFX4 BUFX4_1545 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf2) );
	BUFX4 BUFX4_1546 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf1) );
	BUFX4 BUFX4_1547 ( .gnd(gnd), .vdd(vdd), .A(_14324_), .Y(_14324__bF_buf0) );
	BUFX4 BUFX4_1548 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(_2549__bF_buf4) );
	BUFX4 BUFX4_1549 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(_2549__bF_buf3) );
	BUFX4 BUFX4_1550 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(_2549__bF_buf2) );
	BUFX4 BUFX4_1551 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(_2549__bF_buf1) );
	BUFX4 BUFX4_1552 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(_2549__bF_buf0) );
	BUFX4 BUFX4_1553 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .Y(_2519__bF_buf4) );
	BUFX4 BUFX4_1554 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .Y(_2519__bF_buf3) );
	BUFX4 BUFX4_1555 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .Y(_2519__bF_buf2) );
	BUFX4 BUFX4_1556 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .Y(_2519__bF_buf1) );
	BUFX4 BUFX4_1557 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .Y(_2519__bF_buf0) );
	BUFX4 BUFX4_1558 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_637__bF_buf3) );
	BUFX4 BUFX4_1559 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_637__bF_buf2) );
	BUFX4 BUFX4_1560 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_637__bF_buf1) );
	BUFX4 BUFX4_1561 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_637__bF_buf0) );
	BUFX4 BUFX4_1562 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf5) );
	BUFX4 BUFX4_1563 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf4) );
	BUFX4 BUFX4_1564 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf3) );
	BUFX4 BUFX4_1565 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf2) );
	BUFX4 BUFX4_1566 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf1) );
	BUFX4 BUFX4_1567 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14824__bF_buf0) );
	BUFX4 BUFX4_1568 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9098__bF_buf4) );
	BUFX4 BUFX4_1569 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9098__bF_buf3) );
	BUFX4 BUFX4_1570 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9098__bF_buf2) );
	BUFX4 BUFX4_1571 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9098__bF_buf1) );
	BUFX4 BUFX4_1572 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9098__bF_buf0) );
	BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_), .Y(biu_ins_22_bF_buf3) );
	BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_), .Y(biu_ins_22_bF_buf2) );
	BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_), .Y(biu_ins_22_bF_buf1) );
	BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_), .Y(biu_ins_22_bF_buf0) );
	BUFX4 BUFX4_1573 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11156__bF_buf4) );
	BUFX4 BUFX4_1574 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11156__bF_buf3) );
	BUFX4 BUFX4_1575 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11156__bF_buf2) );
	BUFX4 BUFX4_1576 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11156__bF_buf1) );
	BUFX4 BUFX4_1577 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11156__bF_buf0) );
	BUFX4 BUFX4_1578 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1377__bF_buf3) );
	BUFX4 BUFX4_1579 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1377__bF_buf2) );
	BUFX4 BUFX4_1580 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1377__bF_buf1) );
	BUFX4 BUFX4_1581 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1377__bF_buf0) );
	BUFX4 BUFX4_1582 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .Y(_9105__bF_buf4) );
	BUFX4 BUFX4_1583 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .Y(_9105__bF_buf3) );
	BUFX4 BUFX4_1584 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .Y(_9105__bF_buf2) );
	BUFX4 BUFX4_1585 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .Y(_9105__bF_buf1) );
	BUFX4 BUFX4_1586 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .Y(_9105__bF_buf0) );
	BUFX4 BUFX4_1587 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf5) );
	BUFX4 BUFX4_1588 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf4) );
	BUFX4 BUFX4_1589 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf3) );
	BUFX4 BUFX4_1590 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf2) );
	BUFX4 BUFX4_1591 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf1) );
	BUFX4 BUFX4_1592 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault), .Y(csr_gpr_iu_ins_page_fault_bF_buf0) );
	BUFX4 BUFX4_1593 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .Y(_8192__bF_buf3) );
	BUFX4 BUFX4_1594 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .Y(_8192__bF_buf2) );
	BUFX4 BUFX4_1595 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .Y(_8192__bF_buf1) );
	BUFX4 BUFX4_1596 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .Y(_8192__bF_buf0) );
	BUFX4 BUFX4_1597 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .Y(_8162__bF_buf4) );
	BUFX4 BUFX4_1598 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .Y(_8162__bF_buf3) );
	BUFX4 BUFX4_1599 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .Y(_8162__bF_buf2) );
	BUFX4 BUFX4_1600 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .Y(_8162__bF_buf1) );
	BUFX4 BUFX4_1601 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .Y(_8162__bF_buf0) );
	BUFX4 BUFX4_1602 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf6) );
	BUFX4 BUFX4_1603 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf5) );
	BUFX4 BUFX4_1604 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf4) );
	BUFX4 BUFX4_1605 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf3) );
	BUFX4 BUFX4_1606 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf2) );
	BUFX4 BUFX4_1607 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf1) );
	BUFX4 BUFX4_1608 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7435__bF_buf0) );
	BUFX4 BUFX4_1609 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf14) );
	BUFX4 BUFX4_1610 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf13) );
	BUFX4 BUFX4_1611 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf12) );
	BUFX4 BUFX4_1612 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf11) );
	BUFX4 BUFX4_1613 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf10) );
	BUFX4 BUFX4_1614 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf9) );
	BUFX4 BUFX4_1615 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf8) );
	BUFX4 BUFX4_1616 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf7) );
	BUFX4 BUFX4_1617 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf6) );
	BUFX4 BUFX4_1618 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf5) );
	BUFX4 BUFX4_1619 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf4) );
	BUFX4 BUFX4_1620 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf3) );
	BUFX4 BUFX4_1621 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf2) );
	BUFX4 BUFX4_1622 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf1) );
	BUFX4 BUFX4_1623 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .Y(_7303__bF_buf0) );
	BUFX4 BUFX4_1624 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf6) );
	BUFX4 BUFX4_1625 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf5) );
	BUFX4 BUFX4_1626 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf4) );
	BUFX4 BUFX4_1627 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf3) );
	BUFX4 BUFX4_1628 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf2) );
	BUFX4 BUFX4_1629 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf1) );
	BUFX4 BUFX4_1630 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .Y(_8861__bF_buf0) );
	BUFX4 BUFX4_1631 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf10) );
	BUFX4 BUFX4_1632 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf9) );
	BUFX4 BUFX4_1633 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf8) );
	BUFX4 BUFX4_1634 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf7) );
	BUFX4 BUFX4_1635 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf6) );
	BUFX4 BUFX4_1636 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf5) );
	BUFX4 BUFX4_1637 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf4) );
	BUFX4 BUFX4_1638 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf3) );
	BUFX4 BUFX4_1639 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf2) );
	BUFX4 BUFX4_1640 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf1) );
	BUFX4 BUFX4_1641 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf0) );
	BUFX4 BUFX4_1642 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf15) );
	BUFX4 BUFX4_1643 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf14) );
	BUFX4 BUFX4_1644 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf13) );
	BUFX4 BUFX4_1645 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf12) );
	BUFX4 BUFX4_1646 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf11) );
	BUFX4 BUFX4_1647 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf10) );
	BUFX4 BUFX4_1648 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf9) );
	BUFX4 BUFX4_1649 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf8) );
	BUFX4 BUFX4_1650 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf7) );
	BUFX4 BUFX4_1651 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf6) );
	BUFX4 BUFX4_1652 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf5) );
	BUFX4 BUFX4_1653 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf4) );
	BUFX4 BUFX4_1654 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf3) );
	BUFX4 BUFX4_1655 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf2) );
	BUFX4 BUFX4_1656 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf1) );
	BUFX4 BUFX4_1657 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .Y(_4899__bF_buf0) );
	BUFX4 BUFX4_1658 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .Y(_6492__bF_buf4) );
	BUFX4 BUFX4_1659 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .Y(_6492__bF_buf3) );
	BUFX4 BUFX4_1660 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .Y(_6492__bF_buf2) );
	BUFX4 BUFX4_1661 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .Y(_6492__bF_buf1) );
	BUFX4 BUFX4_1662 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .Y(_6492__bF_buf0) );
	BUFX4 BUFX4_1663 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf5) );
	BUFX4 BUFX4_1664 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf4) );
	BUFX4 BUFX4_1665 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf3) );
	BUFX4 BUFX4_1666 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf2) );
	BUFX4 BUFX4_1667 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf1) );
	BUFX4 BUFX4_1668 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .Y(_7960__bF_buf0) );
	BUFX4 BUFX4_1669 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf5) );
	BUFX4 BUFX4_1670 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf4) );
	BUFX4 BUFX4_1671 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf3) );
	BUFX4 BUFX4_1672 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf2) );
	BUFX4 BUFX4_1673 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf1) );
	BUFX4 BUFX4_1674 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf0) );
	BUFX4 BUFX4_1675 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .Y(_13476__bF_buf3) );
	BUFX4 BUFX4_1676 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .Y(_13476__bF_buf2) );
	BUFX4 BUFX4_1677 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .Y(_13476__bF_buf1) );
	BUFX4 BUFX4_1678 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .Y(_13476__bF_buf0) );
	BUFX4 BUFX4_1679 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf11) );
	BUFX4 BUFX4_1680 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf10) );
	BUFX4 BUFX4_1681 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf9) );
	BUFX4 BUFX4_1682 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf8) );
	BUFX4 BUFX4_1683 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf7) );
	BUFX4 BUFX4_1684 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf6) );
	BUFX4 BUFX4_1685 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf5) );
	BUFX4 BUFX4_1686 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf4) );
	BUFX4 BUFX4_1687 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf3) );
	BUFX4 BUFX4_1688 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf2) );
	BUFX4 BUFX4_1689 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf1) );
	BUFX4 BUFX4_1690 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .Y(_3095__bF_buf0) );
	BUFX4 BUFX4_1691 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .Y(_13416__bF_buf4) );
	BUFX4 BUFX4_1692 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .Y(_13416__bF_buf3) );
	BUFX4 BUFX4_1693 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .Y(_13416__bF_buf2) );
	BUFX4 BUFX4_1694 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .Y(_13416__bF_buf1) );
	BUFX4 BUFX4_1695 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .Y(_13416__bF_buf0) );
	BUFX4 BUFX4_1696 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf6) );
	BUFX4 BUFX4_1697 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf5) );
	BUFX4 BUFX4_1698 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf4) );
	BUFX4 BUFX4_1699 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf3) );
	BUFX4 BUFX4_1700 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf2) );
	BUFX4 BUFX4_1701 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf1) );
	BUFX4 BUFX4_1702 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_), .Y(biu_ins_15_bF_buf0) );
	BUFX4 BUFX4_1703 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_), .Y(addr_csr_17_bF_buf3) );
	BUFX4 BUFX4_1704 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_), .Y(addr_csr_17_bF_buf2) );
	BUFX4 BUFX4_1705 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_), .Y(addr_csr_17_bF_buf1) );
	BUFX4 BUFX4_1706 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_), .Y(addr_csr_17_bF_buf0) );
	BUFX4 BUFX4_1707 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .Y(_11119__bF_buf4) );
	BUFX4 BUFX4_1708 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .Y(_11119__bF_buf3) );
	BUFX4 BUFX4_1709 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .Y(_11119__bF_buf2) );
	BUFX4 BUFX4_1710 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .Y(_11119__bF_buf1) );
	BUFX4 BUFX4_1711 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .Y(_11119__bF_buf0) );
	BUFX4 BUFX4_1712 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf3) );
	BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf2) );
	BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf1) );
	BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf0) );
	BUFX4 BUFX4_1713 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .Y(_2537__bF_buf4) );
	BUFX4 BUFX4_1714 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .Y(_2537__bF_buf3) );
	BUFX4 BUFX4_1715 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .Y(_2537__bF_buf2) );
	BUFX4 BUFX4_1716 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .Y(_2537__bF_buf1) );
	BUFX4 BUFX4_1717 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .Y(_2537__bF_buf0) );
	BUFX4 BUFX4_1718 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .Y(_2507__bF_buf4) );
	BUFX4 BUFX4_1719 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .Y(_2507__bF_buf3) );
	BUFX4 BUFX4_1720 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .Y(_2507__bF_buf2) );
	BUFX4 BUFX4_1721 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .Y(_2507__bF_buf1) );
	BUFX4 BUFX4_1722 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .Y(_2507__bF_buf0) );
	BUFX4 BUFX4_1723 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .Y(_2495__bF_buf4) );
	BUFX4 BUFX4_1724 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .Y(_2495__bF_buf3) );
	BUFX4 BUFX4_1725 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .Y(_2495__bF_buf2) );
	BUFX4 BUFX4_1726 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .Y(_2495__bF_buf1) );
	BUFX4 BUFX4_1727 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .Y(_2495__bF_buf0) );
	BUFX4 BUFX4_1728 ( .gnd(gnd), .vdd(vdd), .A(_854_), .Y(_854__bF_buf4) );
	BUFX4 BUFX4_1729 ( .gnd(gnd), .vdd(vdd), .A(_854_), .Y(_854__bF_buf3) );
	BUFX4 BUFX4_1730 ( .gnd(gnd), .vdd(vdd), .A(_854_), .Y(_854__bF_buf2) );
	BUFX4 BUFX4_1731 ( .gnd(gnd), .vdd(vdd), .A(_854_), .Y(_854__bF_buf1) );
	BUFX4 BUFX4_1732 ( .gnd(gnd), .vdd(vdd), .A(_854_), .Y(_854__bF_buf0) );
	BUFX4 BUFX4_1733 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .Y(_13441__bF_buf4) );
	BUFX4 BUFX4_1734 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .Y(_13441__bF_buf3) );
	BUFX4 BUFX4_1735 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .Y(_13441__bF_buf2) );
	BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .Y(_13441__bF_buf1) );
	BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .Y(_13441__bF_buf0) );
	BUFX4 BUFX4_1736 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .Y(_4931__bF_buf4) );
	BUFX4 BUFX4_1737 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .Y(_4931__bF_buf3) );
	BUFX4 BUFX4_1738 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .Y(_4931__bF_buf2) );
	BUFX4 BUFX4_1739 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .Y(_4931__bF_buf1) );
	BUFX4 BUFX4_1740 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .Y(_4931__bF_buf0) );
	BUFX4 BUFX4_1741 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf8) );
	BUFX4 BUFX4_1742 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf7) );
	BUFX4 BUFX4_1743 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf6) );
	BUFX4 BUFX4_1744 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf5) );
	BUFX4 BUFX4_1745 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf4) );
	BUFX4 BUFX4_1746 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf3) );
	BUFX4 BUFX4_1747 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf2) );
	BUFX4 BUFX4_1748 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf1) );
	BUFX4 BUFX4_1749 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .Y(_2995__bF_buf0) );
	BUFX4 BUFX4_1750 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf7) );
	BUFX4 BUFX4_1751 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf6) );
	BUFX4 BUFX4_1752 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf5) );
	BUFX4 BUFX4_1753 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf4) );
	BUFX4 BUFX4_1754 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf3) );
	BUFX4 BUFX4_1755 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf2) );
	BUFX4 BUFX4_1756 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf1) );
	BUFX4 BUFX4_1757 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .Y(_2694__bF_buf0) );
	BUFX4 BUFX4_1758 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf4) );
	BUFX4 BUFX4_1759 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf3) );
	BUFX4 BUFX4_1760 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf2) );
	BUFX4 BUFX4_1761 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf1) );
	BUFX4 BUFX4_1762 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf0) );
	BUFX4 BUFX4_1763 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_), .Y(biu_exce_chk_statu_biu_4_bF_buf3) );
	BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_), .Y(biu_exce_chk_statu_biu_4_bF_buf2) );
	BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_), .Y(biu_exce_chk_statu_biu_4_bF_buf1) );
	BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_), .Y(biu_exce_chk_statu_biu_4_bF_buf0) );
	BUFX4 BUFX4_1764 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf5) );
	BUFX4 BUFX4_1765 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf4) );
	BUFX4 BUFX4_1766 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf3) );
	BUFX4 BUFX4_1767 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf2) );
	BUFX4 BUFX4_1768 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf1) );
	BUFX4 BUFX4_1769 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .Y(_1004__bF_buf0) );
	BUFX4 BUFX4_1770 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .Y(_8486__bF_buf3) );
	BUFX4 BUFX4_1771 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .Y(_8486__bF_buf2) );
	BUFX4 BUFX4_1772 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .Y(_8486__bF_buf1) );
	BUFX4 BUFX4_1773 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .Y(_8486__bF_buf0) );
	BUFX4 BUFX4_1774 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf8) );
	BUFX4 BUFX4_1775 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf7) );
	BUFX4 BUFX4_1776 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf6) );
	BUFX4 BUFX4_1777 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf5) );
	BUFX4 BUFX4_1778 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf4) );
	BUFX4 BUFX4_1779 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf3) );
	BUFX4 BUFX4_1780 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf2) );
	BUFX4 BUFX4_1781 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf1) );
	BUFX4 BUFX4_1782 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .Y(_7428__bF_buf0) );
	BUFX4 BUFX4_1783 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6159__bF_buf4) );
	BUFX4 BUFX4_1784 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6159__bF_buf3) );
	BUFX4 BUFX4_1785 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6159__bF_buf2) );
	BUFX4 BUFX4_1786 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6159__bF_buf1) );
	BUFX4 BUFX4_1787 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6159__bF_buf0) );
	BUFX4 BUFX4_1788 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .Y(_2460__bF_buf4) );
	BUFX4 BUFX4_1789 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .Y(_2460__bF_buf3) );
	BUFX4 BUFX4_1790 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .Y(_2460__bF_buf2) );
	BUFX4 BUFX4_1791 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .Y(_2460__bF_buf1) );
	BUFX4 BUFX4_1792 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .Y(_2460__bF_buf0) );
	BUFX4 BUFX4_1793 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2731__bF_buf4) );
	BUFX4 BUFX4_1794 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2731__bF_buf3) );
	BUFX4 BUFX4_1795 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2731__bF_buf2) );
	BUFX4 BUFX4_1796 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2731__bF_buf1) );
	BUFX4 BUFX4_1797 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2731__bF_buf0) );
	BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf3) );
	BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf2) );
	BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf1) );
	BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf0) );
	BUFX4 BUFX4_1798 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .Y(_9021__bF_buf4) );
	BUFX4 BUFX4_1799 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .Y(_9021__bF_buf3) );
	BUFX4 BUFX4_1800 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .Y(_9021__bF_buf2) );
	BUFX4 BUFX4_1801 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .Y(_9021__bF_buf1) );
	BUFX4 BUFX4_1802 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .Y(_9021__bF_buf0) );
	BUFX4 BUFX4_1803 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .Y(_6226__bF_buf4) );
	BUFX4 BUFX4_1804 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .Y(_6226__bF_buf3) );
	BUFX4 BUFX4_1805 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .Y(_6226__bF_buf2) );
	BUFX4 BUFX4_1806 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .Y(_6226__bF_buf1) );
	BUFX4 BUFX4_1807 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .Y(_6226__bF_buf0) );
	BUFX4 BUFX4_1808 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .Y(_6425__bF_buf4) );
	BUFX4 BUFX4_1809 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .Y(_6425__bF_buf3) );
	BUFX4 BUFX4_1810 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .Y(_6425__bF_buf2) );
	BUFX4 BUFX4_1811 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .Y(_6425__bF_buf1) );
	BUFX4 BUFX4_1812 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .Y(_6425__bF_buf0) );
	BUFX4 BUFX4_1813 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .Y(_13397__bF_buf4) );
	BUFX4 BUFX4_1814 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .Y(_13397__bF_buf3) );
	BUFX4 BUFX4_1815 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .Y(_13397__bF_buf2) );
	BUFX4 BUFX4_1816 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .Y(_13397__bF_buf1) );
	BUFX4 BUFX4_1817 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .Y(_13397__bF_buf0) );
	BUFX4 BUFX4_1818 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .Y(_12297__bF_buf4) );
	BUFX4 BUFX4_1819 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .Y(_12297__bF_buf3) );
	BUFX4 BUFX4_1820 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .Y(_12297__bF_buf2) );
	BUFX4 BUFX4_1821 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .Y(_12297__bF_buf1) );
	BUFX4 BUFX4_1822 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .Y(_12297__bF_buf0) );
	BUFX4 BUFX4_1823 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf5) );
	BUFX4 BUFX4_1824 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf4) );
	BUFX4 BUFX4_1825 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf3) );
	BUFX4 BUFX4_1826 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf2) );
	BUFX4 BUFX4_1827 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf1) );
	BUFX4 BUFX4_1828 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .Y(_9019__bF_buf0) );
	BUFX4 BUFX4_1829 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .Y(_13464__bF_buf3) );
	BUFX4 BUFX4_1830 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .Y(_13464__bF_buf2) );
	BUFX4 BUFX4_1831 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .Y(_13464__bF_buf1) );
	BUFX4 BUFX4_1832 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .Y(_13464__bF_buf0) );
	BUFX4 BUFX4_1833 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf7) );
	BUFX4 BUFX4_1834 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf6) );
	BUFX4 BUFX4_1835 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf5) );
	BUFX4 BUFX4_1836 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf4) );
	BUFX4 BUFX4_1837 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf3) );
	BUFX4 BUFX4_1838 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf2) );
	BUFX4 BUFX4_1839 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf1) );
	BUFX4 BUFX4_1840 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .Y(_13392__bF_buf0) );
	BUFX4 BUFX4_1841 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(_2525__bF_buf4) );
	BUFX4 BUFX4_1842 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(_2525__bF_buf3) );
	BUFX4 BUFX4_1843 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(_2525__bF_buf2) );
	BUFX4 BUFX4_1844 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(_2525__bF_buf1) );
	BUFX4 BUFX4_1845 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(_2525__bF_buf0) );
	BUFX4 BUFX4_1846 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf5) );
	BUFX4 BUFX4_1847 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf4) );
	BUFX4 BUFX4_1848 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf3) );
	BUFX4 BUFX4_1849 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf2) );
	BUFX4 BUFX4_1850 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf1) );
	BUFX4 BUFX4_1851 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .Y(_8419__bF_buf0) );
	BUFX4 BUFX4_1852 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf5) );
	BUFX4 BUFX4_1853 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf4) );
	BUFX4 BUFX4_1854 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf3) );
	BUFX4 BUFX4_1855 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf2) );
	BUFX4 BUFX4_1856 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf1) );
	BUFX4 BUFX4_1857 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .Y(_8118__bF_buf0) );
	BUFX4 BUFX4_1858 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2483__bF_buf4) );
	BUFX4 BUFX4_1859 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2483__bF_buf3) );
	BUFX4 BUFX4_1860 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2483__bF_buf2) );
	BUFX4 BUFX4_1861 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2483__bF_buf1) );
	BUFX4 BUFX4_1862 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2483__bF_buf0) );
	BUFX4 BUFX4_1863 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf6) );
	BUFX4 BUFX4_1864 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf5) );
	BUFX4 BUFX4_1865 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf4) );
	BUFX4 BUFX4_1866 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf3) );
	BUFX4 BUFX4_1867 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf2) );
	BUFX4 BUFX4_1868 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf1) );
	BUFX4 BUFX4_1869 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_8618__bF_buf0) );
	BUFX4 BUFX4_1870 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .Y(_7319__bF_buf4) );
	BUFX4 BUFX4_1871 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .Y(_7319__bF_buf3) );
	BUFX4 BUFX4_1872 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .Y(_7319__bF_buf2) );
	BUFX4 BUFX4_1873 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .Y(_7319__bF_buf1) );
	BUFX4 BUFX4_1874 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .Y(_7319__bF_buf0) );
	BUFX4 BUFX4_1875 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .Y(_9273__bF_buf3) );
	BUFX4 BUFX4_1876 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .Y(_9273__bF_buf2) );
	BUFX4 BUFX4_1877 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .Y(_9273__bF_buf1) );
	BUFX4 BUFX4_1878 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .Y(_9273__bF_buf0) );
	BUFX4 BUFX4_1879 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf7) );
	BUFX4 BUFX4_1880 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf6) );
	BUFX4 BUFX4_1881 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf5) );
	BUFX4 BUFX4_1882 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf4) );
	BUFX4 BUFX4_1883 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf3) );
	BUFX4 BUFX4_1884 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf2) );
	BUFX4 BUFX4_1885 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf1) );
	BUFX4 BUFX4_1886 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .Y(_8847__bF_buf0) );
	BUFX4 BUFX4_1887 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf7) );
	BUFX4 BUFX4_1888 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf6) );
	BUFX4 BUFX4_1889 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf5) );
	BUFX4 BUFX4_1890 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf4) );
	BUFX4 BUFX4_1891 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf3) );
	BUFX4 BUFX4_1892 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf2) );
	BUFX4 BUFX4_1893 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf1) );
	BUFX4 BUFX4_1894 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_710__bF_buf0) );
	BUFX4 BUFX4_1895 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .Y(_8516__bF_buf3) );
	BUFX4 BUFX4_1896 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .Y(_8516__bF_buf2) );
	BUFX4 BUFX4_1897 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .Y(_8516__bF_buf1) );
	BUFX4 BUFX4_1898 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .Y(_8516__bF_buf0) );
	BUFX4 BUFX4_1899 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_), .Y(csr_gpr_iu_csr_priv_d_1_bF_buf3) );
	BUFX4 BUFX4_1900 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_), .Y(csr_gpr_iu_csr_priv_d_1_bF_buf2) );
	BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_), .Y(csr_gpr_iu_csr_priv_d_1_bF_buf1) );
	BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_), .Y(csr_gpr_iu_csr_priv_d_1_bF_buf0) );
	BUFX4 BUFX4_1901 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .Y(_1221__bF_buf4) );
	BUFX4 BUFX4_1902 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .Y(_1221__bF_buf3) );
	BUFX4 BUFX4_1903 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .Y(_1221__bF_buf2) );
	BUFX4 BUFX4_1904 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .Y(_1221__bF_buf1) );
	BUFX4 BUFX4_1905 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .Y(_1221__bF_buf0) );
	BUFX4 BUFX4_1906 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf6) );
	BUFX4 BUFX4_1907 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf5) );
	BUFX4 BUFX4_1908 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf4) );
	BUFX4 BUFX4_1909 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf3) );
	BUFX4 BUFX4_1910 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf2) );
	BUFX4 BUFX4_1911 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf1) );
	BUFX4 BUFX4_1912 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .Y(_8372__bF_buf0) );
	BUFX4 BUFX4_1913 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf5) );
	BUFX4 BUFX4_1914 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf4) );
	BUFX4 BUFX4_1915 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf3) );
	BUFX4 BUFX4_1916 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf2) );
	BUFX4 BUFX4_1917 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf1) );
	BUFX4 BUFX4_1918 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .Y(_14328__bF_buf0) );
	BUFX4 BUFX4_1919 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_), .Y(biu_ins_26_bF_buf3) );
	BUFX4 BUFX4_1920 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_), .Y(biu_ins_26_bF_buf2) );
	BUFX4 BUFX4_1921 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_), .Y(biu_ins_26_bF_buf1) );
	BUFX4 BUFX4_1922 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_), .Y(biu_ins_26_bF_buf0) );
	BUFX4 BUFX4_1923 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf6) );
	BUFX4 BUFX4_1924 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf5) );
	BUFX4 BUFX4_1925 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf4) );
	BUFX4 BUFX4_1926 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf3) );
	BUFX4 BUFX4_1927 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf2) );
	BUFX4 BUFX4_1928 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf1) );
	BUFX4 BUFX4_1929 ( .gnd(gnd), .vdd(vdd), .A(addi), .Y(addi_bF_buf0) );
	BUFX4 BUFX4_1930 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .Y(_14323__bF_buf3) );
	BUFX4 BUFX4_1931 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .Y(_14323__bF_buf2) );
	BUFX4 BUFX4_1932 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .Y(_14323__bF_buf1) );
	BUFX4 BUFX4_1933 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .Y(_14323__bF_buf0) );
	BUFX4 BUFX4_1934 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .Y(_12086__bF_buf3) );
	BUFX4 BUFX4_1935 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .Y(_12086__bF_buf2) );
	BUFX4 BUFX4_1936 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .Y(_12086__bF_buf1) );
	BUFX4 BUFX4_1937 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .Y(_12086__bF_buf0) );
	BUFX4 BUFX4_1938 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_666__bF_buf4) );
	BUFX4 BUFX4_1939 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_666__bF_buf3) );
	BUFX4 BUFX4_1940 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_666__bF_buf2) );
	BUFX4 BUFX4_1941 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_666__bF_buf1) );
	BUFX4 BUFX4_1942 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_666__bF_buf0) );
	BUFX4 BUFX4_1943 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .Y(_1249__bF_buf3) );
	BUFX4 BUFX4_1944 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .Y(_1249__bF_buf2) );
	BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .Y(_1249__bF_buf1) );
	BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .Y(_1249__bF_buf0) );
	BUFX4 BUFX4_1945 ( .gnd(gnd), .vdd(vdd), .A(addp), .Y(addp_bF_buf4) );
	BUFX4 BUFX4_1946 ( .gnd(gnd), .vdd(vdd), .A(addp), .Y(addp_bF_buf3) );
	BUFX4 BUFX4_1947 ( .gnd(gnd), .vdd(vdd), .A(addp), .Y(addp_bF_buf2) );
	BUFX4 BUFX4_1948 ( .gnd(gnd), .vdd(vdd), .A(addp), .Y(addp_bF_buf1) );
	BUFX4 BUFX4_1949 ( .gnd(gnd), .vdd(vdd), .A(addp), .Y(addp_bF_buf0) );
	BUFX4 BUFX4_1950 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf15) );
	BUFX4 BUFX4_1951 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf14) );
	BUFX4 BUFX4_1952 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf13) );
	BUFX4 BUFX4_1953 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf12) );
	BUFX4 BUFX4_1954 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf11) );
	BUFX4 BUFX4_1955 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf10) );
	BUFX4 BUFX4_1956 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf9) );
	BUFX4 BUFX4_1957 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf8) );
	BUFX4 BUFX4_1958 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf7) );
	BUFX4 BUFX4_1959 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf6) );
	BUFX4 BUFX4_1960 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf5) );
	BUFX4 BUFX4_1961 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf4) );
	BUFX4 BUFX4_1962 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf3) );
	BUFX4 BUFX4_1963 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf2) );
	BUFX4 BUFX4_1964 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf1) );
	BUFX4 BUFX4_1965 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .Y(_3113__bF_buf0) );
	BUFX4 BUFX4_1966 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_835__bF_buf4) );
	BUFX4 BUFX4_1967 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_835__bF_buf3) );
	BUFX4 BUFX4_1968 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_835__bF_buf2) );
	BUFX4 BUFX4_1969 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_835__bF_buf1) );
	BUFX4 BUFX4_1970 ( .gnd(gnd), .vdd(vdd), .A(_835_), .Y(_835__bF_buf0) );
	BUFX4 BUFX4_1971 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_), .Y(biu_ins_21_bF_buf3) );
	BUFX4 BUFX4_1972 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_), .Y(biu_ins_21_bF_buf2) );
	BUFX4 BUFX4_1973 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_), .Y(biu_ins_21_bF_buf1) );
	BUFX4 BUFX4_1974 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_), .Y(biu_ins_21_bF_buf0) );
	BUFX4 BUFX4_1975 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_), .Y(addr_csr_23_bF_buf3) );
	BUFX4 BUFX4_1976 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_), .Y(addr_csr_23_bF_buf2) );
	BUFX4 BUFX4_1977 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_), .Y(addr_csr_23_bF_buf1) );
	BUFX4 BUFX4_1978 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_), .Y(addr_csr_23_bF_buf0) );
	BUFX4 BUFX4_1979 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2543__bF_buf4) );
	BUFX4 BUFX4_1980 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2543__bF_buf3) );
	BUFX4 BUFX4_1981 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2543__bF_buf2) );
	BUFX4 BUFX4_1982 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2543__bF_buf1) );
	BUFX4 BUFX4_1983 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2543__bF_buf0) );
	BUFX4 BUFX4_1984 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf4) );
	BUFX4 BUFX4_1985 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf3) );
	BUFX4 BUFX4_1986 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf2) );
	BUFX4 BUFX4_1987 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf1) );
	BUFX4 BUFX4_1988 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf0) );
	BUFX4 BUFX4_1989 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .Y(_7439__bF_buf4) );
	BUFX4 BUFX4_1990 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .Y(_7439__bF_buf3) );
	BUFX4 BUFX4_1991 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .Y(_7439__bF_buf2) );
	BUFX4 BUFX4_1992 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .Y(_7439__bF_buf1) );
	BUFX4 BUFX4_1993 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .Y(_7439__bF_buf0) );
	BUFX4 BUFX4_1994 ( .gnd(gnd), .vdd(vdd), .A(_10182_), .Y(_10182__bF_buf3) );
	BUFX4 BUFX4_1995 ( .gnd(gnd), .vdd(vdd), .A(_10182_), .Y(_10182__bF_buf2) );
	BUFX4 BUFX4_1996 ( .gnd(gnd), .vdd(vdd), .A(_10182_), .Y(_10182__bF_buf1) );
	BUFX4 BUFX4_1997 ( .gnd(gnd), .vdd(vdd), .A(_10182_), .Y(_10182__bF_buf0) );
	BUFX4 BUFX4_1998 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf5) );
	BUFX4 BUFX4_1999 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf4) );
	BUFX4 BUFX4_2000 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf3) );
	BUFX4 BUFX4_2001 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf2) );
	BUFX4 BUFX4_2002 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf1) );
	BUFX4 BUFX4_2003 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .Y(_8233__bF_buf0) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(data_rd_0_), .Y(_0_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_0_), .Y(_1_) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .Y(_2_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(biu_exce_chk_opc_2_), .Y(_3_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lb), .B(csr_gpr_iu_ins_dec_lh), .Y(_4_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf3), .B(_4_), .C(_3_), .Y(_5_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .Y(_6_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(_6_), .Y(_7_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(csr_gpr_iu_ins_dec_lb), .Y(_8_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_7_), .Y(_9_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(csr_gpr_iu_ins_dec_lh), .C(_3_), .Y(_10_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_5_), .C(_9_), .Y(_11_) );
	MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_0_), .S(_11_), .Y(csr_gpr_iu_data_gpr_0_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(data_rd_1_), .Y(_12_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_1_), .Y(_13_) );
	MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_12_), .S(_11_), .Y(csr_gpr_iu_data_gpr_1_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(data_rd_2_), .Y(_14_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_2_), .Y(_15_) );
	MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_14_), .S(_11_), .Y(csr_gpr_iu_data_gpr_2_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(data_rd_3_), .Y(_16_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .Y(_17_) );
	MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_16_), .S(_11_), .Y(csr_gpr_iu_data_gpr_3_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(data_rd_4_), .Y(_18_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .Y(_19_) );
	MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_18_), .S(_11_), .Y(csr_gpr_iu_data_gpr_4_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(data_rd_5_), .Y(_20_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_5_), .Y(_21_) );
	MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_20_), .S(_11_), .Y(csr_gpr_iu_data_gpr_5_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(data_rd_6_), .Y(_22_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_6_), .Y(_23_) );
	MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_22_), .S(_11_), .Y(csr_gpr_iu_data_gpr_6_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(data_rd_7_), .Y(_24_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .Y(_25_) );
	MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_24_), .S(_11_), .Y(csr_gpr_iu_data_gpr_7_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .Y(_26_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(biu_exce_chk_opc_2_), .Y(_27_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(_27__bF_buf3), .Y(_28_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .B(csr_gpr_iu_ins_dec_lb), .Y(_29_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(_2__bF_buf2), .C(_29_), .Y(_30_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_30__bF_buf3), .B(biu_biu_data_out_7_bF_buf2), .C(_28__bF_buf3), .Y(_31_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(biu_exce_chk_opc_0_), .C(biu_exce_chk_opc_2_), .Y(_32_) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_32__bF_buf3), .Y(_33_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lb), .Y(_34_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_8_), .C(_34_), .D(_28__bF_buf2), .Y(_35_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(data_rd_8_), .B(_33_), .C(_35__bF_buf3), .Y(_36_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_3_), .C(_31_), .D(_36_), .Y(csr_gpr_iu_data_gpr_8_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_9_), .Y(_37_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(data_rd_9_), .B(_33_), .C(_35__bF_buf2), .Y(_38_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_3_), .C(_31_), .D(_38_), .Y(csr_gpr_iu_data_gpr_9_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_10_), .Y(_39_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(data_rd_10_), .B(_33_), .C(_35__bF_buf1), .Y(_40_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_3_), .C(_31_), .D(_40_), .Y(csr_gpr_iu_data_gpr_10_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_11_), .Y(_41_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(data_rd_11_), .B(_33_), .C(_35__bF_buf0), .Y(_42_) );
	AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_3_), .C(_31_), .D(_42_), .Y(csr_gpr_iu_data_gpr_11_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_12_), .Y(_43_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(data_rd_12_), .B(_33_), .C(_35__bF_buf3), .Y(_44_) );
	AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_3_), .C(_31_), .D(_44_), .Y(csr_gpr_iu_data_gpr_12_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_13_), .Y(_45_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(data_rd_13_), .B(_33_), .C(_35__bF_buf2), .Y(_46_) );
	AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_3_), .C(_31_), .D(_46_), .Y(csr_gpr_iu_data_gpr_13_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_14_), .Y(_47_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(data_rd_14_), .B(_33_), .C(_35__bF_buf1), .Y(_48_) );
	AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_3_), .C(_31_), .D(_48_), .Y(csr_gpr_iu_data_gpr_14_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .Y(_49_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(data_rd_15_), .B(_33_), .C(_35__bF_buf0), .Y(_50_) );
	AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_3_), .C(_31_), .D(_50_), .Y(csr_gpr_iu_data_gpr_15_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lh), .B(biu_biu_data_out_15_), .C(_28__bF_buf1), .Y(_51_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_16_), .Y(_52_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf1), .B(_27__bF_buf2), .C(data_rd_16_), .Y(_53_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_32__bF_buf2), .C(_53_), .Y(_54_) );
	AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf1), .B(_30__bF_buf2), .C(_54_), .D(_35__bF_buf3), .Y(_55_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf0), .B(_55_), .C(_51_), .Y(csr_gpr_iu_data_gpr_16_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_17_), .Y(_56_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf0), .B(_27__bF_buf1), .C(data_rd_17_), .Y(_57_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_32__bF_buf1), .C(_57_), .Y(_58_) );
	AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf0), .B(_30__bF_buf1), .C(_58_), .D(_35__bF_buf2), .Y(_59_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf3), .B(_59_), .C(_51_), .Y(csr_gpr_iu_data_gpr_17_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_18_), .Y(_60_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf3), .B(_27__bF_buf0), .C(data_rd_18_), .Y(_61_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_32__bF_buf0), .C(_61_), .Y(_62_) );
	AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .B(_30__bF_buf0), .C(_62_), .D(_35__bF_buf1), .Y(_63_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf2), .B(_63_), .C(_51_), .Y(csr_gpr_iu_data_gpr_18_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_19_), .Y(_64_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf2), .B(_27__bF_buf3), .C(data_rd_19_), .Y(_65_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_32__bF_buf3), .C(_65_), .Y(_66_) );
	AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf2), .B(_30__bF_buf3), .C(_66_), .D(_35__bF_buf0), .Y(_67_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf1), .B(_67_), .C(_51_), .Y(csr_gpr_iu_data_gpr_19_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_20_), .Y(_68_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf1), .B(_27__bF_buf2), .C(data_rd_20_), .Y(_69_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_32__bF_buf2), .C(_69_), .Y(_70_) );
	AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf1), .B(_30__bF_buf2), .C(_70_), .D(_35__bF_buf3), .Y(_71_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf0), .B(_71_), .C(_51_), .Y(csr_gpr_iu_data_gpr_20_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_21_), .Y(_72_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf0), .B(_27__bF_buf1), .C(data_rd_21_), .Y(_73_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_32__bF_buf1), .C(_73_), .Y(_74_) );
	AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf0), .B(_30__bF_buf1), .C(_74_), .D(_35__bF_buf2), .Y(_75_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf3), .B(_75_), .C(_51_), .Y(csr_gpr_iu_data_gpr_21_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_22_), .Y(_76_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf3), .B(_27__bF_buf0), .C(data_rd_22_), .Y(_77_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_32__bF_buf0), .C(_77_), .Y(_78_) );
	AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .B(_30__bF_buf0), .C(_78_), .D(_35__bF_buf1), .Y(_79_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf2), .B(_79_), .C(_51_), .Y(csr_gpr_iu_data_gpr_22_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_23_), .Y(_80_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf2), .B(_27__bF_buf3), .C(data_rd_23_), .Y(_81_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_32__bF_buf3), .C(_81_), .Y(_82_) );
	AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf2), .B(_30__bF_buf3), .C(_82_), .D(_35__bF_buf0), .Y(_83_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf1), .B(_83_), .C(_51_), .Y(csr_gpr_iu_data_gpr_23_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_24_), .Y(_84_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf1), .B(_27__bF_buf2), .C(data_rd_24_), .Y(_85_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_32__bF_buf2), .C(_85_), .Y(_86_) );
	AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf1), .B(_30__bF_buf2), .C(_86_), .D(_35__bF_buf3), .Y(_87_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf0), .B(_87_), .C(_51_), .Y(csr_gpr_iu_data_gpr_24_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_25_), .Y(_88_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf0), .B(_27__bF_buf1), .C(data_rd_25_), .Y(_89_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_32__bF_buf1), .C(_89_), .Y(_90_) );
	AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf0), .B(_30__bF_buf1), .C(_90_), .D(_35__bF_buf2), .Y(_91_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf3), .B(_91_), .C(_51_), .Y(csr_gpr_iu_data_gpr_25_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_26_), .Y(_92_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf3), .B(_27__bF_buf0), .C(data_rd_26_), .Y(_93_) );
	OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_32__bF_buf0), .C(_93_), .Y(_94_) );
	AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .B(_30__bF_buf0), .C(_94_), .D(_35__bF_buf1), .Y(_95_) );
	OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf2), .B(_95_), .C(_51_), .Y(csr_gpr_iu_data_gpr_26_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_27_), .Y(_96_) );
	OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf2), .B(_27__bF_buf3), .C(data_rd_27_), .Y(_97_) );
	OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_32__bF_buf3), .C(_97_), .Y(_98_) );
	AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf2), .B(_30__bF_buf3), .C(_98_), .D(_35__bF_buf0), .Y(_99_) );
	OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf1), .B(_99_), .C(_51_), .Y(csr_gpr_iu_data_gpr_27_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_28_), .Y(_100_) );
	OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf1), .B(_27__bF_buf2), .C(data_rd_28_), .Y(_101_) );
	OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_32__bF_buf2), .C(_101_), .Y(_102_) );
	AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf1), .B(_30__bF_buf2), .C(_102_), .D(_35__bF_buf3), .Y(_103_) );
	OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf0), .B(_103_), .C(_51_), .Y(csr_gpr_iu_data_gpr_28_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_29_), .Y(_104_) );
	OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf0), .B(_27__bF_buf1), .C(data_rd_29_), .Y(_105_) );
	OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_32__bF_buf1), .C(_105_), .Y(_106_) );
	AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf0), .B(_30__bF_buf1), .C(_106_), .D(_35__bF_buf2), .Y(_107_) );
	OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf3), .B(_107_), .C(_51_), .Y(csr_gpr_iu_data_gpr_29_) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_30_), .Y(_108_) );
	OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf3), .B(_27__bF_buf0), .C(data_rd_30_), .Y(_109_) );
	OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_32__bF_buf0), .C(_109_), .Y(_110_) );
	AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .B(_30__bF_buf0), .C(_110_), .D(_35__bF_buf1), .Y(_111_) );
	OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf2), .B(_111_), .C(_51_), .Y(csr_gpr_iu_data_gpr_30_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_31_), .Y(_112_) );
	OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2__bF_buf2), .B(_27__bF_buf3), .C(data_rd_31_), .Y(_113_) );
	OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_32__bF_buf3), .C(_113_), .Y(_114_) );
	AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf2), .B(_30__bF_buf3), .C(_114_), .D(_35__bF_buf0), .Y(_115_) );
	OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_28__bF_buf1), .B(_115_), .C(_51_), .Y(csr_gpr_iu_data_gpr_31_) );
	BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(_116__0_), .Y(haddr[0]) );
	BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(_116__1_), .Y(haddr[1]) );
	BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(_116__2_), .Y(haddr[2]) );
	BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(_116__3_), .Y(haddr[3]) );
	BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(_116__4_), .Y(haddr[4]) );
	BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(_116__5_), .Y(haddr[5]) );
	BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(_116__6_), .Y(haddr[6]) );
	BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(_116__7_), .Y(haddr[7]) );
	BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(_116__8_), .Y(haddr[8]) );
	BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(_116__9_), .Y(haddr[9]) );
	BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(_116__10_), .Y(haddr[10]) );
	BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(_116__11_), .Y(haddr[11]) );
	BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(_116__12_), .Y(haddr[12]) );
	BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(_116__13_), .Y(haddr[13]) );
	BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(_116__14_), .Y(haddr[14]) );
	BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(_116__15_), .Y(haddr[15]) );
	BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(_116__16_), .Y(haddr[16]) );
	BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(_116__17_), .Y(haddr[17]) );
	BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(_116__18_), .Y(haddr[18]) );
	BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(_116__19_), .Y(haddr[19]) );
	BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(_116__20_), .Y(haddr[20]) );
	BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(_116__21_), .Y(haddr[21]) );
	BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(_116__22_), .Y(haddr[22]) );
	BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(_116__23_), .Y(haddr[23]) );
	BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(_116__24_), .Y(haddr[24]) );
	BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(_116__25_), .Y(haddr[25]) );
	BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(_116__26_), .Y(haddr[26]) );
	BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(_116__27_), .Y(haddr[27]) );
	BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(_116__28_), .Y(haddr[28]) );
	BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(_116__29_), .Y(haddr[29]) );
	BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(_116__30_), .Y(haddr[30]) );
	BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(_116__31_), .Y(haddr[31]) );
	BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(_116__32_), .Y(haddr[32]) );
	BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(_116__33_), .Y(haddr[33]) );
	BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hburst[0]) );
	BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hburst[1]) );
	BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hburst[2]) );
	BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hmastlock) );
	BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(hprot[0]) );
	BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(hprot[1]) );
	BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hprot[2]) );
	BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hprot[3]) );
	BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(_117__0_), .Y(hsize[0]) );
	BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(_117__1_), .Y(hsize[1]) );
	BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(htrans[0]) );
	BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(_118__1_), .Y(htrans[1]) );
	BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(_119__0_), .Y(hwdata[0]) );
	BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(_119__1_), .Y(hwdata[1]) );
	BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(_119__2_), .Y(hwdata[2]) );
	BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(_119__3_), .Y(hwdata[3]) );
	BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(_119__4_), .Y(hwdata[4]) );
	BUFX2 BUFX2_173 ( .gnd(gnd), .vdd(vdd), .A(_119__5_), .Y(hwdata[5]) );
	BUFX2 BUFX2_174 ( .gnd(gnd), .vdd(vdd), .A(_119__6_), .Y(hwdata[6]) );
	BUFX2 BUFX2_175 ( .gnd(gnd), .vdd(vdd), .A(_119__7_), .Y(hwdata[7]) );
	BUFX2 BUFX2_176 ( .gnd(gnd), .vdd(vdd), .A(_119__8_), .Y(hwdata[8]) );
	BUFX2 BUFX2_177 ( .gnd(gnd), .vdd(vdd), .A(_119__9_), .Y(hwdata[9]) );
	BUFX2 BUFX2_178 ( .gnd(gnd), .vdd(vdd), .A(_119__10_), .Y(hwdata[10]) );
	BUFX2 BUFX2_179 ( .gnd(gnd), .vdd(vdd), .A(_119__11_), .Y(hwdata[11]) );
	BUFX2 BUFX2_180 ( .gnd(gnd), .vdd(vdd), .A(_119__12_), .Y(hwdata[12]) );
	BUFX2 BUFX2_181 ( .gnd(gnd), .vdd(vdd), .A(_119__13_), .Y(hwdata[13]) );
	BUFX2 BUFX2_182 ( .gnd(gnd), .vdd(vdd), .A(_119__14_), .Y(hwdata[14]) );
	BUFX2 BUFX2_183 ( .gnd(gnd), .vdd(vdd), .A(_119__15_), .Y(hwdata[15]) );
	BUFX2 BUFX2_184 ( .gnd(gnd), .vdd(vdd), .A(_119__16_), .Y(hwdata[16]) );
	BUFX2 BUFX2_185 ( .gnd(gnd), .vdd(vdd), .A(_119__17_), .Y(hwdata[17]) );
	BUFX2 BUFX2_186 ( .gnd(gnd), .vdd(vdd), .A(_119__18_), .Y(hwdata[18]) );
	BUFX2 BUFX2_187 ( .gnd(gnd), .vdd(vdd), .A(_119__19_), .Y(hwdata[19]) );
	BUFX2 BUFX2_188 ( .gnd(gnd), .vdd(vdd), .A(_119__20_), .Y(hwdata[20]) );
	BUFX2 BUFX2_189 ( .gnd(gnd), .vdd(vdd), .A(_119__21_), .Y(hwdata[21]) );
	BUFX2 BUFX2_190 ( .gnd(gnd), .vdd(vdd), .A(_119__22_), .Y(hwdata[22]) );
	BUFX2 BUFX2_191 ( .gnd(gnd), .vdd(vdd), .A(_119__23_), .Y(hwdata[23]) );
	BUFX2 BUFX2_192 ( .gnd(gnd), .vdd(vdd), .A(_119__24_), .Y(hwdata[24]) );
	BUFX2 BUFX2_193 ( .gnd(gnd), .vdd(vdd), .A(_119__25_), .Y(hwdata[25]) );
	BUFX2 BUFX2_194 ( .gnd(gnd), .vdd(vdd), .A(_119__26_), .Y(hwdata[26]) );
	BUFX2 BUFX2_195 ( .gnd(gnd), .vdd(vdd), .A(_119__27_), .Y(hwdata[27]) );
	BUFX2 BUFX2_196 ( .gnd(gnd), .vdd(vdd), .A(_119__28_), .Y(hwdata[28]) );
	BUFX2 BUFX2_197 ( .gnd(gnd), .vdd(vdd), .A(_119__29_), .Y(hwdata[29]) );
	BUFX2 BUFX2_198 ( .gnd(gnd), .vdd(vdd), .A(_119__30_), .Y(hwdata[30]) );
	BUFX2 BUFX2_199 ( .gnd(gnd), .vdd(vdd), .A(_119__31_), .Y(hwdata[31]) );
	BUFX2 BUFX2_200 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(hwrite) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .Y(_628_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .Y(_629_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .B(biu_exce_chk_statu_biu_2_), .Y(_630_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_630_), .Y(_631_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_631_), .Y(_632_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_632_), .Y(_633_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf3), .Y(_634_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .Y(_635_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_635_), .Y(_636_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf3), .B(_636_), .Y(_637_) );
	INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf3), .Y(_638_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_633_), .Y(biu_rdy_biu) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(biu_exce_chk_statu_biu_1_), .Y(_639_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_639_), .Y(_640_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .Y(_641_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(biu_exce_chk_statu_biu_2_), .Y(_642_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_642_), .Y(_643_) );
	INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(_643_), .Y(_644_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_644_), .Y(_645_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf6), .Y(_646_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf2), .B(_635_), .Y(_647_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_648_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf2), .B(_648_), .Y(_649_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_649_), .Y(_650_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf1), .B(_634_), .Y(_651_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(_651_), .Y(_652_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_652_), .Y(_653_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_653_), .Y(_654_) );
	INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf0), .Y(_655_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(_634_), .Y(_656_) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_656_), .Y(_657_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_657_), .Y(_658_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_636_), .Y(_659_) );
	OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_658_), .C(_643_), .Y(_660_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_654_), .C(_660_), .Y(_661_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf3), .B(_657_), .Y(_662_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_648_), .Y(_663_) );
	OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .C(_643_), .Y(_664_) );
	OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_638_), .C(_664_), .Y(_665_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_661_), .Y(_666_) );
	INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_666__bF_buf4), .Y(_667_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .Y(_668_) );
	OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_661_), .C(_668_), .Y(_669_) );
	OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_1_), .B(_667_), .C(_669_), .Y(_670_) );
	OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_644_), .C(_670_), .Y(_671_) );
	OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .B(_646_), .C(_671_), .Y(_672_) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_672_), .Y(_116__1_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .Y(_673_) );
	OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_661_), .C(_673_), .Y(_674_) );
	OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_0_), .B(_667_), .C(_674_), .Y(_675_) );
	OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_644_), .C(_675_), .Y(_676_) );
	OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .B(_646_), .C(_676_), .Y(_677_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_677_), .Y(_116__0_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(biu_exce_chk_statu_cpu_1_), .Y(_678_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(biu_exce_chk_statu_cpu_3_), .Y(_679_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .Y(_680_) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .Y(_681_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_681_), .Y(_682_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .C(_682_), .Y(_683_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_673_), .Y(_684_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(biu_exce_chk_opc_1_), .Y(_685_) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .Y(_686_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(_686_), .Y(_687_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(addr_csr_0_), .Y(_688_) );
	AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_685_), .C(_688_), .D(_687_), .Y(_689_) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .Y(_690_) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .Y(_691_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(_691_), .Y(_692_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_692_), .Y(_693_) );
	OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_689_), .C(_683_), .Y(biu_addr_mis) );
	INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_633_), .Y(_694_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(_632_), .Y(_695_) );
	INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(_695_), .Y(_696_) );
	OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_694_), .C(_662_), .Y(_697_) );
	INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_662_), .Y(_698_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_639_), .Y(_699_) );
	OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_699_), .C(_646_), .Y(_700_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(_641_), .Y(_701_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_640_), .Y(_702_) );
	INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(_702_), .Y(_703_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(_631_), .Y(_704_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(_704_), .Y(_705_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_698_), .Y(_706_) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_706_), .Y(_707_) );
	OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_703_), .C(_707_), .Y(_708_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_708_), .Y(_709_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_697_), .Y(_710_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_710__bF_buf7), .Y(_711_) );
	OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_710__bF_buf6), .C(_711_), .Y(biu_addr_mmu_in_0_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_710__bF_buf5), .Y(_712_) );
	OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_710__bF_buf4), .C(_712_), .Y(biu_addr_mmu_in_1_) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .Y(_713_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_710__bF_buf3), .Y(_714_) );
	OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_710__bF_buf2), .C(_714_), .Y(biu_addr_mmu_in_2_) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .Y(_715_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_710__bF_buf1), .Y(_716_) );
	OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_710__bF_buf0), .C(_716_), .Y(biu_addr_mmu_in_3_) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .Y(_717_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_710__bF_buf7), .Y(_718_) );
	OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_710__bF_buf6), .C(_718_), .Y(biu_addr_mmu_in_4_) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .Y(_719_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_710__bF_buf5), .Y(_720_) );
	OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_710__bF_buf4), .C(_720_), .Y(biu_addr_mmu_in_5_) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .Y(_721_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_710__bF_buf3), .Y(_722_) );
	OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_710__bF_buf2), .C(_722_), .Y(biu_addr_mmu_in_6_) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .Y(_723_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_710__bF_buf1), .Y(_724_) );
	OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_710__bF_buf0), .C(_724_), .Y(biu_addr_mmu_in_7_) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .Y(_725_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_710__bF_buf7), .Y(_726_) );
	OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_710__bF_buf6), .C(_726_), .Y(biu_addr_mmu_in_8_) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .Y(_727_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_710__bF_buf5), .Y(_728_) );
	OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_710__bF_buf4), .C(_728_), .Y(biu_addr_mmu_in_9_) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .Y(_729_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_710__bF_buf3), .Y(_730_) );
	OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_710__bF_buf2), .C(_730_), .Y(biu_addr_mmu_in_10_) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .Y(_731_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .B(_710__bF_buf1), .Y(_732_) );
	OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_710__bF_buf0), .C(_732_), .Y(biu_addr_mmu_in_11_) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .Y(_733_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_710__bF_buf7), .Y(_734_) );
	OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_710__bF_buf6), .C(_734_), .Y(biu_addr_mmu_in_12_) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .Y(_735_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_710__bF_buf5), .Y(_736_) );
	OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_710__bF_buf4), .C(_736_), .Y(biu_addr_mmu_in_13_) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .Y(_737_) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_710__bF_buf3), .Y(_738_) );
	OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_710__bF_buf2), .C(_738_), .Y(biu_addr_mmu_in_14_) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .Y(_739_) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf3), .B(_710__bF_buf1), .Y(_740_) );
	OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_710__bF_buf0), .C(_740_), .Y(biu_addr_mmu_in_15_) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .Y(_741_) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_710__bF_buf7), .Y(_742_) );
	OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_710__bF_buf6), .C(_742_), .Y(biu_addr_mmu_in_16_) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .Y(_743_) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf3), .B(_710__bF_buf5), .Y(_744_) );
	OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_710__bF_buf4), .C(_744_), .Y(biu_addr_mmu_in_17_) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .Y(_745_) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_710__bF_buf3), .Y(_746_) );
	OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_710__bF_buf2), .C(_746_), .Y(biu_addr_mmu_in_18_) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .Y(_747_) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_710__bF_buf1), .Y(_748_) );
	OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_710__bF_buf0), .C(_748_), .Y(biu_addr_mmu_in_19_) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .Y(_749_) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_710__bF_buf7), .Y(_750_) );
	OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_710__bF_buf6), .C(_750_), .Y(biu_addr_mmu_in_20_) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .Y(_751_) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_710__bF_buf5), .Y(_752_) );
	OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_710__bF_buf4), .C(_752_), .Y(biu_addr_mmu_in_21_) );
	INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .Y(_753_) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_710__bF_buf3), .Y(_754_) );
	OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_710__bF_buf2), .C(_754_), .Y(biu_addr_mmu_in_22_) );
	INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .Y(_755_) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf3), .B(_710__bF_buf1), .Y(_756_) );
	OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_710__bF_buf0), .C(_756_), .Y(biu_addr_mmu_in_23_) );
	INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .Y(_757_) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_710__bF_buf7), .Y(_758_) );
	OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_710__bF_buf6), .C(_758_), .Y(biu_addr_mmu_in_24_) );
	INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .Y(_759_) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_710__bF_buf5), .Y(_760_) );
	OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_710__bF_buf4), .C(_760_), .Y(biu_addr_mmu_in_25_) );
	INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .Y(_761_) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .B(_710__bF_buf3), .Y(_762_) );
	OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_710__bF_buf2), .C(_762_), .Y(biu_addr_mmu_in_26_) );
	INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .Y(_763_) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_710__bF_buf1), .Y(_764_) );
	OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_710__bF_buf0), .C(_764_), .Y(biu_addr_mmu_in_27_) );
	INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .Y(_765_) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_710__bF_buf7), .Y(_766_) );
	OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_710__bF_buf6), .C(_766_), .Y(biu_addr_mmu_in_28_) );
	INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .Y(_767_) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_710__bF_buf5), .Y(_768_) );
	OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_710__bF_buf4), .C(_768_), .Y(biu_addr_mmu_in_29_) );
	INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .Y(_769_) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_710__bF_buf3), .Y(_770_) );
	OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_710__bF_buf2), .C(_770_), .Y(biu_addr_mmu_in_30_) );
	INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .Y(_771_) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf3), .B(_710__bF_buf1), .Y(_772_) );
	OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_710__bF_buf0), .C(_772_), .Y(biu_addr_mmu_in_31_) );
	MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_2_), .B(addr_csr_2_), .S(_666__bF_buf3), .Y(_773_) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(_645__bF_buf5), .Y(_774_) );
	OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf4), .B(_773_), .C(_774_), .Y(_116__2_) );
	MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_3_), .B(addr_csr_3_), .S(_666__bF_buf2), .Y(_775_) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .B(_645__bF_buf3), .Y(_776_) );
	OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf2), .B(_775_), .C(_776_), .Y(_116__3_) );
	MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_4_), .B(addr_csr_4_), .S(_666__bF_buf1), .Y(_777_) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .B(_645__bF_buf1), .Y(_778_) );
	OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf0), .B(_777_), .C(_778_), .Y(_116__4_) );
	MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_5_), .B(addr_csr_5_), .S(_666__bF_buf0), .Y(_779_) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .B(_645__bF_buf6), .Y(_780_) );
	OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf5), .B(_779_), .C(_780_), .Y(_116__5_) );
	MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_6_), .B(addr_csr_6_), .S(_666__bF_buf4), .Y(_781_) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .B(_645__bF_buf4), .Y(_782_) );
	OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf3), .B(_781_), .C(_782_), .Y(_116__6_) );
	MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_7_), .B(addr_csr_7_), .S(_666__bF_buf3), .Y(_783_) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .B(_645__bF_buf2), .Y(_784_) );
	OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf1), .B(_783_), .C(_784_), .Y(_116__7_) );
	MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_8_), .B(addr_csr_8_), .S(_666__bF_buf2), .Y(_785_) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .B(_645__bF_buf0), .Y(_786_) );
	OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf6), .B(_785_), .C(_786_), .Y(_116__8_) );
	MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_9_), .B(addr_csr_9_), .S(_666__bF_buf1), .Y(_787_) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .B(_645__bF_buf5), .Y(_788_) );
	OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf4), .B(_787_), .C(_788_), .Y(_116__9_) );
	MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_10_), .B(addr_csr_10_), .S(_666__bF_buf0), .Y(_789_) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(_645__bF_buf3), .Y(_790_) );
	OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf2), .B(_789_), .C(_790_), .Y(_116__10_) );
	MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_11_), .B(addr_csr_11_), .S(_666__bF_buf4), .Y(_791_) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(_645__bF_buf1), .Y(_792_) );
	OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf0), .B(_791_), .C(_792_), .Y(_116__11_) );
	MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_12_), .B(addr_csr_12_), .S(_666__bF_buf3), .Y(_793_) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .B(_645__bF_buf6), .Y(_794_) );
	OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf5), .B(_793_), .C(_794_), .Y(_116__12_) );
	MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_13_), .B(addr_csr_13_bF_buf2), .S(_666__bF_buf2), .Y(_795_) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(_645__bF_buf4), .Y(_796_) );
	OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf3), .B(_795_), .C(_796_), .Y(_116__13_) );
	MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_14_), .B(addr_csr_14_), .S(_666__bF_buf1), .Y(_797_) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(_645__bF_buf2), .Y(_798_) );
	OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf1), .B(_797_), .C(_798_), .Y(_116__14_) );
	MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_15_), .B(addr_csr_15_bF_buf2), .S(_666__bF_buf0), .Y(_799_) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .B(_645__bF_buf0), .Y(_800_) );
	OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf6), .B(_799_), .C(_800_), .Y(_116__15_) );
	MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_16_), .B(addr_csr_16_), .S(_666__bF_buf4), .Y(_801_) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .B(_645__bF_buf5), .Y(_802_) );
	OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf4), .B(_801_), .C(_802_), .Y(_116__16_) );
	MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_17_), .B(addr_csr_17_bF_buf2), .S(_666__bF_buf3), .Y(_803_) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(_645__bF_buf3), .Y(_804_) );
	OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf2), .B(_803_), .C(_804_), .Y(_116__17_) );
	MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_18_), .B(addr_csr_18_), .S(_666__bF_buf2), .Y(_805_) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(_645__bF_buf1), .Y(_806_) );
	OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf0), .B(_805_), .C(_806_), .Y(_116__18_) );
	MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_19_), .B(addr_csr_19_bF_buf2), .S(_666__bF_buf1), .Y(_807_) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .B(_645__bF_buf6), .Y(_808_) );
	OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf5), .B(_807_), .C(_808_), .Y(_116__19_) );
	MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_20_), .B(addr_csr_20_), .S(_666__bF_buf0), .Y(_809_) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_645__bF_buf4), .Y(_810_) );
	OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf3), .B(_809_), .C(_810_), .Y(_116__20_) );
	MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_21_), .B(addr_csr_21_bF_buf2), .S(_666__bF_buf4), .Y(_811_) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .B(_645__bF_buf2), .Y(_812_) );
	OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf1), .B(_811_), .C(_812_), .Y(_116__21_) );
	MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_22_), .B(addr_csr_22_), .S(_666__bF_buf3), .Y(_813_) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_645__bF_buf0), .Y(_814_) );
	OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf6), .B(_813_), .C(_814_), .Y(_116__22_) );
	MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_23_), .B(addr_csr_23_bF_buf2), .S(_666__bF_buf2), .Y(_815_) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .B(_645__bF_buf5), .Y(_816_) );
	OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf4), .B(_815_), .C(_816_), .Y(_116__23_) );
	MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_24_), .B(addr_csr_24_), .S(_666__bF_buf1), .Y(_817_) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .B(_645__bF_buf3), .Y(_818_) );
	OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf2), .B(_817_), .C(_818_), .Y(_116__24_) );
	MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_25_), .B(addr_csr_25_bF_buf2), .S(_666__bF_buf0), .Y(_819_) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .B(_645__bF_buf1), .Y(_820_) );
	OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf0), .B(_819_), .C(_820_), .Y(_116__25_) );
	MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_26_), .B(addr_csr_26_), .S(_666__bF_buf4), .Y(_821_) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(_645__bF_buf6), .Y(_822_) );
	OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf5), .B(_821_), .C(_822_), .Y(_116__26_) );
	MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_27_), .B(addr_csr_27_bF_buf2), .S(_666__bF_buf3), .Y(_823_) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .B(_645__bF_buf4), .Y(_824_) );
	OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf3), .B(_823_), .C(_824_), .Y(_116__27_) );
	MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_28_), .B(addr_csr_28_), .S(_666__bF_buf2), .Y(_825_) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .B(_645__bF_buf2), .Y(_826_) );
	OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf1), .B(_825_), .C(_826_), .Y(_116__28_) );
	MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_29_), .B(addr_csr_29_bF_buf2), .S(_666__bF_buf1), .Y(_827_) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(_645__bF_buf0), .Y(_828_) );
	OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf6), .B(_827_), .C(_828_), .Y(_116__29_) );
	MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_30_), .B(addr_csr_30_), .S(_666__bF_buf0), .Y(_829_) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(_645__bF_buf5), .Y(_830_) );
	OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf4), .B(_829_), .C(_830_), .Y(_116__30_) );
	MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_31_), .B(addr_csr_31_bF_buf2), .S(_666__bF_buf4), .Y(_831_) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .B(_645__bF_buf3), .Y(_832_) );
	OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf2), .B(_831_), .C(_832_), .Y(_116__31_) );
	OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_644_), .C(biu_addr_mmu_32_), .Y(_833_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_667_), .Y(_116__32_) );
	OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_644_), .C(biu_addr_mmu_33_), .Y(_834_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_667_), .Y(_116__33_) );
	OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf2), .B(_636_), .C(_632_), .Y(_835_) );
	INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_0_), .Y(_836_) );
	INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_632_), .Y(_837_) );
	OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf2), .B(_837__bF_buf3), .C(_836_), .Y(_838_) );
	OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_0_), .B(_835__bF_buf4), .C(_838_), .Y(_839_) );
	INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_663_), .Y(_840_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_840_), .Y(_841_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_635_), .Y(_842_) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf1), .B(_842_), .Y(_843_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_703_), .Y(_844_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_841_), .Y(_845_) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_643_), .Y(_846_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_846_), .Y(_847_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_840_), .Y(_848_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_848_), .Y(_849_) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_849_), .Y(_850_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_116__1_), .Y(_851_) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_851_), .Y(_852_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_116__0_), .Y(_853_) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_853_), .Y(_854_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_677_), .Y(_855_) );
	OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_844_), .C(_855_), .Y(_856_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf3), .B(_852_), .C(_854__bF_buf4), .Y(_857_) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_857_), .Y(biu_ahb_data_in_0_) );
	INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_1_), .Y(_858_) );
	OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf1), .B(_837__bF_buf2), .C(_858_), .Y(_859_) );
	OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_1_), .B(_835__bF_buf3), .C(_859_), .Y(_860_) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_857_), .Y(biu_ahb_data_in_1_) );
	INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_2_), .Y(_861_) );
	OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf0), .B(_837__bF_buf1), .C(_861_), .Y(_862_) );
	OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_2_), .B(_835__bF_buf2), .C(_862_), .Y(_863_) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_857_), .Y(biu_ahb_data_in_2_) );
	INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_3_), .Y(_864_) );
	OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf3), .B(_837__bF_buf0), .C(_864_), .Y(_865_) );
	OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_3_), .B(_835__bF_buf1), .C(_865_), .Y(_866_) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_857_), .Y(biu_ahb_data_in_3_) );
	INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_4_), .Y(_867_) );
	OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf2), .B(_837__bF_buf3), .C(_867_), .Y(_868_) );
	OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_4_), .B(_835__bF_buf0), .C(_868_), .Y(_869_) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_857_), .Y(biu_ahb_data_in_4_) );
	INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_5_), .Y(_870_) );
	OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf1), .B(_837__bF_buf2), .C(_870_), .Y(_871_) );
	OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_5_), .B(_835__bF_buf4), .C(_871_), .Y(_872_) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_857_), .Y(biu_ahb_data_in_5_) );
	MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_6_), .B(biu_mmu_pte_new_7_bF_buf4), .S(_835__bF_buf3), .Y(_873_) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_857_), .Y(biu_ahb_data_in_6_) );
	INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_7_), .Y(_874_) );
	OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf0), .B(_837__bF_buf1), .C(_874_), .Y(_875_) );
	OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(_835__bF_buf2), .C(_875_), .Y(_876_) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_857_), .Y(biu_ahb_data_in_7_) );
	INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_8_), .Y(_877_) );
	OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf3), .B(_837__bF_buf0), .C(_877_), .Y(_878_) );
	OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_8_), .B(_835__bF_buf1), .C(_878_), .Y(_879_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_852_), .C(_879_), .D(_857_), .Y(biu_ahb_data_in_8_) );
	INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_9_), .Y(_880_) );
	OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf2), .B(_837__bF_buf3), .C(_880_), .Y(_881_) );
	OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_9_), .B(_835__bF_buf0), .C(_881_), .Y(_882_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_860_), .C(_882_), .D(_857_), .Y(biu_ahb_data_in_9_) );
	INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_10_), .Y(_883_) );
	OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf1), .B(_837__bF_buf2), .C(_883_), .Y(_884_) );
	OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_10_), .B(_835__bF_buf4), .C(_884_), .Y(_885_) );
	OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_863_), .C(_885_), .D(_857_), .Y(biu_ahb_data_in_10_) );
	INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_11_), .Y(_886_) );
	OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf0), .B(_837__bF_buf1), .C(_886_), .Y(_887_) );
	OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_11_), .B(_835__bF_buf3), .C(_887_), .Y(_888_) );
	OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_866_), .C(_888_), .D(_857_), .Y(biu_ahb_data_in_11_) );
	INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_12_), .Y(_889_) );
	OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf3), .B(_837__bF_buf0), .C(_889_), .Y(_890_) );
	OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_12_), .B(_835__bF_buf2), .C(_890_), .Y(_891_) );
	OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_869_), .C(_891_), .D(_857_), .Y(biu_ahb_data_in_12_) );
	INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_13_), .Y(_892_) );
	OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf2), .B(_837__bF_buf3), .C(_892_), .Y(_893_) );
	OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_13_), .B(_835__bF_buf1), .C(_893_), .Y(_894_) );
	OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_872_), .C(_894_), .D(_857_), .Y(biu_ahb_data_in_13_) );
	INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_14_), .Y(_895_) );
	OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf1), .B(_837__bF_buf2), .C(_895_), .Y(_896_) );
	OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_14_), .B(_835__bF_buf0), .C(_896_), .Y(_897_) );
	OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_873_), .C(_897_), .D(_857_), .Y(biu_ahb_data_in_14_) );
	INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_15_), .Y(_898_) );
	OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf0), .B(_837__bF_buf1), .C(_898_), .Y(_899_) );
	OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_15_), .B(_835__bF_buf4), .C(_899_), .Y(_900_) );
	OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_876_), .C(_900_), .D(_857_), .Y(biu_ahb_data_in_15_) );
	INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_852_), .Y(_901_) );
	INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_839_), .Y(_902_) );
	INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf2), .Y(_903_) );
	MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_16_), .B(biu_mmu_pte_new_16_), .S(_835__bF_buf3), .Y(_904_) );
	OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_903_), .C(_854__bF_buf3), .Y(_905_) );
	OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_854__bF_buf2), .C(_905_), .Y(_906_) );
	INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_907_) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_901_), .Y(_908_) );
	OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_906_), .C(_908_), .Y(biu_ahb_data_in_16_) );
	INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_860_), .Y(_909_) );
	MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_17_), .B(biu_mmu_pte_new_17_), .S(_835__bF_buf2), .Y(_910_) );
	OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_903_), .C(_854__bF_buf1), .Y(_911_) );
	OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf0), .B(_909_), .C(_911_), .Y(_912_) );
	INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_882_), .Y(_913_) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_913_), .B(_901_), .Y(_914_) );
	OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_912_), .C(_914_), .Y(biu_ahb_data_in_17_) );
	INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_863_), .Y(_915_) );
	MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_18_), .B(biu_mmu_pte_new_18_), .S(_835__bF_buf1), .Y(_916_) );
	OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_903_), .C(_854__bF_buf4), .Y(_917_) );
	OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf3), .B(_915_), .C(_917_), .Y(_918_) );
	INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_885_), .Y(_919_) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_901_), .Y(_920_) );
	OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_918_), .C(_920_), .Y(biu_ahb_data_in_18_) );
	INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_866_), .Y(_921_) );
	MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_19_), .B(biu_mmu_pte_new_19_), .S(_835__bF_buf0), .Y(_922_) );
	OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_903_), .C(_854__bF_buf2), .Y(_923_) );
	OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf1), .B(_921_), .C(_923_), .Y(_924_) );
	INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_925_) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_901_), .Y(_926_) );
	OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_924_), .C(_926_), .Y(biu_ahb_data_in_19_) );
	INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_869_), .Y(_927_) );
	MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_20_), .B(biu_mmu_pte_new_20_), .S(_835__bF_buf4), .Y(_928_) );
	OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_903_), .C(_854__bF_buf0), .Y(_929_) );
	OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf4), .B(_927_), .C(_929_), .Y(_930_) );
	INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_891_), .Y(_931_) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_901_), .Y(_932_) );
	OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_930_), .C(_932_), .Y(biu_ahb_data_in_20_) );
	INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_872_), .Y(_933_) );
	MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_21_), .B(biu_mmu_pte_new_21_), .S(_835__bF_buf3), .Y(_934_) );
	OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_903_), .C(_854__bF_buf3), .Y(_935_) );
	OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf2), .B(_933_), .C(_935_), .Y(_936_) );
	INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_894_), .Y(_937_) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_901_), .Y(_938_) );
	OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_936_), .C(_938_), .Y(biu_ahb_data_in_21_) );
	NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_854__bF_buf1), .Y(_939_) );
	OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_637__bF_buf3), .B(_837__bF_buf0), .C(biu_biu_data_in_22_), .Y(_940_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_22_), .B(_632_), .C(_638_), .Y(_941_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_941_), .C(_903_), .Y(_942_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_854__bF_buf0), .C(_939_), .Y(_943_) );
	INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_897_), .Y(_944_) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_901_), .Y(_945_) );
	OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_943_), .C(_945_), .Y(biu_ahb_data_in_22_) );
	INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_946_) );
	MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_23_), .B(biu_mmu_pte_new_23_), .S(_835__bF_buf2), .Y(_947_) );
	OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_903_), .C(_854__bF_buf4), .Y(_948_) );
	OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf3), .B(_946_), .C(_948_), .Y(_949_) );
	INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_950_) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_901_), .Y(_951_) );
	OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_949_), .C(_951_), .Y(biu_ahb_data_in_23_) );
	NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_116__1_), .B(_116__0_), .Y(_952_) );
	OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf1), .B(biu_exce_chk_statu_biu_5_), .C(_632_), .Y(_953_) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_694_), .Y(_954_) );
	INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_658_), .Y(_955_) );
	INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_659_), .Y(_956_) );
	NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_644_), .Y(_957_) );
	INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_957_), .Y(_958_) );
	OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_703_), .C(_958_), .Y(_959_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_696_), .C(_959_), .Y(_960_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(_954_), .C(_960_), .Y(_961_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_850_), .C(_961_), .Y(_962_) );
	MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_24_), .B(biu_mmu_pte_new_24_), .S(_835__bF_buf1), .Y(_963_) );
	INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_963_), .Y(_964_) );
	OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_856__bF_buf1), .C(_854__bF_buf2), .Y(_965_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf0), .B(_964_), .C(_965_), .Y(_966_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_852_), .Y(_967_) );
	OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf1), .B(_907_), .C(_967_), .Y(_968_) );
	OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_963_), .C(_966_), .D(_968_), .Y(biu_ahb_data_in_24_) );
	MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_25_), .B(biu_mmu_pte_new_25_), .S(_835__bF_buf0), .Y(_969_) );
	INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_969_), .Y(_970_) );
	OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_856__bF_buf3), .C(_854__bF_buf0), .Y(_971_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf2), .B(_970_), .C(_971_), .Y(_972_) );
	OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf4), .B(_913_), .C(_967_), .Y(_973_) );
	OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_969_), .C(_972_), .D(_973_), .Y(biu_ahb_data_in_25_) );
	MUX2X1 MUX2X1_49 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_26_), .B(biu_mmu_pte_new_26_), .S(_835__bF_buf4), .Y(_974_) );
	INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_974_), .Y(_975_) );
	OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_856__bF_buf1), .C(_854__bF_buf3), .Y(_976_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf0), .B(_975_), .C(_976_), .Y(_977_) );
	OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf2), .B(_919_), .C(_967_), .Y(_978_) );
	OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_974_), .C(_977_), .D(_978_), .Y(biu_ahb_data_in_26_) );
	MUX2X1 MUX2X1_50 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_27_), .B(biu_mmu_pte_new_27_), .S(_835__bF_buf3), .Y(_979_) );
	INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_979_), .Y(_980_) );
	OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_856__bF_buf3), .C(_854__bF_buf1), .Y(_981_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf2), .B(_980_), .C(_981_), .Y(_982_) );
	OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf0), .B(_925_), .C(_967_), .Y(_983_) );
	OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_979_), .C(_982_), .D(_983_), .Y(biu_ahb_data_in_27_) );
	MUX2X1 MUX2X1_51 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_28_), .B(biu_mmu_pte_new_28_), .S(_835__bF_buf2), .Y(_984_) );
	INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_984_), .Y(_985_) );
	OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_856__bF_buf1), .C(_854__bF_buf4), .Y(_986_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf0), .B(_985_), .C(_986_), .Y(_987_) );
	OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf3), .B(_931_), .C(_967_), .Y(_988_) );
	OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_984_), .C(_987_), .D(_988_), .Y(biu_ahb_data_in_28_) );
	MUX2X1 MUX2X1_52 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_29_), .B(biu_mmu_pte_new_29_), .S(_835__bF_buf1), .Y(_989_) );
	INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_989_), .Y(_990_) );
	OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_856__bF_buf3), .C(_854__bF_buf2), .Y(_991_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf2), .B(_990_), .C(_991_), .Y(_992_) );
	OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf1), .B(_937_), .C(_967_), .Y(_993_) );
	OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_989_), .C(_992_), .D(_993_), .Y(biu_ahb_data_in_29_) );
	MUX2X1 MUX2X1_53 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_30_), .B(biu_mmu_pte_new_30_), .S(_835__bF_buf0), .Y(_994_) );
	INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_994_), .Y(_995_) );
	OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_856__bF_buf1), .C(_854__bF_buf0), .Y(_996_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf0), .B(_995_), .C(_996_), .Y(_997_) );
	OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf4), .B(_944_), .C(_967_), .Y(_998_) );
	OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_994_), .C(_997_), .D(_998_), .Y(biu_ahb_data_in_30_) );
	MUX2X1 MUX2X1_54 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_31_), .B(biu_mmu_pte_new_31_), .S(_835__bF_buf4), .Y(_999_) );
	INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_1000_) );
	OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_856__bF_buf3), .C(_854__bF_buf3), .Y(_1001_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_856__bF_buf2), .B(_1000_), .C(_1001_), .Y(_1002_) );
	OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_854__bF_buf2), .B(_950_), .C(_967_), .Y(_1003_) );
	OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_999_), .C(_1002_), .D(_1003_), .Y(biu_ahb_data_in_31_) );
	NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(biu_rdy_biu), .Y(_1004_) );
	NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_0_), .B(_1004__bF_buf5), .Y(_1005_) );
	NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .B(_687_), .Y(_1006_) );
	INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .Y(_1007_) );
	NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_851_), .Y(_1008_) );
	INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .Y(_1009_) );
	INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_16_), .Y(_1010_) );
	NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_853_), .Y(_1011_) );
	INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .Y(_1012_) );
	NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(_1012_), .Y(_1013_) );
	NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .B(_1013_), .Y(_1014_) );
	INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .Y(_1015_) );
	NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_853_), .Y(_1016_) );
	NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1016_), .Y(_1017_) );
	INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(_855_), .Y(_1018_) );
	NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .Y(_1019_) );
	MUX2X1 MUX2X1_55 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_24_), .B(biu_ahb_data_out_0_), .S(_1019_), .Y(_1020_) );
	NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_851_), .Y(_1021_) );
	INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1022_) );
	NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_1017_), .Y(_1023_) );
	AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1017_), .C(_1023_), .D(_1020_), .Y(_1024_) );
	INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_8_), .Y(_1025_) );
	OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_1015_), .C(_851_), .Y(_1026_) );
	INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .Y(_1027_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_1025_), .C(_1004__bF_buf4), .Y(_1028_) );
	OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf3), .B(_1024_), .C(_1028_), .Y(_1029_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_1005_), .C(rst_bF_buf70), .Y(_121__0_) );
	NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_1_), .B(_1004__bF_buf3), .Y(_1030_) );
	INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(_1004__bF_buf2), .Y(_1031_) );
	INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_9_), .Y(_1032_) );
	INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_25_), .Y(_1033_) );
	INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1034_) );
	OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .C(biu_ahb_data_out_1_), .Y(_1035_) );
	OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_1034_), .C(_1035_), .Y(_1036_) );
	AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_17_), .B(_1017_), .C(_1023_), .D(_1036_), .Y(_1037_) );
	OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_1026_), .C(_1009__bF_buf2), .D(_1037_), .Y(_1038_) );
	NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf3), .B(_1038_), .Y(_1039_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1030_), .C(rst_bF_buf69), .Y(_121__1_) );
	NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_2_), .B(_1004__bF_buf1), .Y(_1040_) );
	INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_10_), .Y(_1041_) );
	INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_26_), .Y(_1042_) );
	OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .C(biu_ahb_data_out_2_), .Y(_1043_) );
	OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1034_), .C(_1043_), .Y(_1044_) );
	AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_18_), .B(_1017_), .C(_1023_), .D(_1044_), .Y(_1045_) );
	OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_1026_), .C(_1009__bF_buf1), .D(_1045_), .Y(_1046_) );
	NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(_1046_), .Y(_1047_) );
	AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .B(_1040_), .C(rst_bF_buf68), .Y(_121__2_) );
	NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .B(_1004__bF_buf0), .Y(_1048_) );
	INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_11_), .Y(_1049_) );
	INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_27_), .Y(_1050_) );
	OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .C(biu_ahb_data_out_3_), .Y(_1051_) );
	OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1034_), .C(_1051_), .Y(_1052_) );
	AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_19_), .B(_1017_), .C(_1023_), .D(_1052_), .Y(_1053_) );
	OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1026_), .C(_1009__bF_buf0), .D(_1053_), .Y(_1054_) );
	NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf1), .B(_1054_), .Y(_1055_) );
	AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1048_), .C(rst_bF_buf67), .Y(_121__3_) );
	NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .B(_1004__bF_buf5), .Y(_1056_) );
	INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_12_), .Y(_1057_) );
	INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_28_), .Y(_1058_) );
	OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .C(biu_ahb_data_out_4_), .Y(_1059_) );
	OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1034_), .C(_1059_), .Y(_1060_) );
	AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_20_), .B(_1017_), .C(_1023_), .D(_1060_), .Y(_1061_) );
	OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1026_), .C(_1009__bF_buf3), .D(_1061_), .Y(_1062_) );
	NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf0), .B(_1062_), .Y(_1063_) );
	AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1056_), .C(rst_bF_buf66), .Y(_121__4_) );
	NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_5_), .B(_1004__bF_buf4), .Y(_1064_) );
	INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_13_), .Y(_124_) );
	INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_29_), .Y(_125_) );
	OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1018_), .C(biu_ahb_data_out_5_), .Y(_126_) );
	OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_1034_), .C(_126_), .Y(_127_) );
	AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_21_), .B(_1017_), .C(_1023_), .D(_127_), .Y(_128_) );
	OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_1026_), .C(_1009__bF_buf2), .D(_128_), .Y(_129_) );
	NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf3), .B(_129_), .Y(_130_) );
	AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_1064_), .C(rst_bF_buf65), .Y(_121__5_) );
	NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_6_), .B(_1004__bF_buf3), .Y(_131_) );
	INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_22_), .Y(_132_) );
	MUX2X1 MUX2X1_56 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_30_), .B(biu_ahb_data_out_6_), .S(_1019_), .Y(_133_) );
	AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_1017_), .C(_1023_), .D(_133_), .Y(_134_) );
	INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_14_), .Y(_135_) );
	AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_135_), .C(_1004__bF_buf2), .Y(_136_) );
	OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf1), .B(_134_), .C(_136_), .Y(_137_) );
	AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_131_), .C(rst_bF_buf64), .Y(_121__6_) );
	NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf1), .B(_1004__bF_buf1), .Y(_138_) );
	INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_23_), .Y(_139_) );
	MUX2X1 MUX2X1_57 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_31_), .B(biu_ahb_data_out_7_), .S(_1019_), .Y(_140_) );
	AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_1017_), .C(_1023_), .D(_140_), .Y(_141_) );
	INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_15_), .Y(_142_) );
	AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_142_), .C(_1004__bF_buf0), .Y(_143_) );
	OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf0), .B(_141_), .C(_143_), .Y(_144_) );
	AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_138_), .C(rst_bF_buf63), .Y(_121__7_) );
	NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .B(_1004__bF_buf5), .Y(_145_) );
	OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1014_), .C(_1023_), .Y(_146_) );
	INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .Y(_147_) );
	AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_24_), .C(_1009__bF_buf3), .Y(_148_) );
	OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_146_), .C(_148_), .Y(_149_) );
	AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_1031__bF_buf2), .Y(_150_) );
	OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_16_), .B(_1008_), .C(_150_), .Y(_151_) );
	AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_145_), .C(rst_bF_buf62), .Y(_121__8_) );
	NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_9_), .B(_1004__bF_buf4), .Y(_152_) );
	AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_25_), .C(_1009__bF_buf2), .Y(_153_) );
	OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_146_), .C(_153_), .Y(_154_) );
	AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf1), .B(biu_ahb_data_out_17_), .Y(_155_) );
	NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1004__bF_buf3), .B(_1009__bF_buf1), .Y(_156_) );
	OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .C(_154_), .Y(_157_) );
	AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_152_), .C(rst_bF_buf61), .Y(_121__9_) );
	NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_10_), .B(_1004__bF_buf2), .Y(_158_) );
	AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_26_), .C(_1009__bF_buf0), .Y(_159_) );
	OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_146_), .C(_159_), .Y(_160_) );
	AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf0), .B(biu_ahb_data_out_18_), .Y(_161_) );
	OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_161_), .C(_160_), .Y(_162_) );
	AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_158_), .C(rst_bF_buf60), .Y(_121__10_) );
	NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_11_), .B(_1004__bF_buf1), .Y(_163_) );
	AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_27_), .C(_1009__bF_buf3), .Y(_164_) );
	OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_146_), .C(_164_), .Y(_165_) );
	AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf3), .B(biu_ahb_data_out_19_), .Y(_166_) );
	OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_166_), .C(_165_), .Y(_167_) );
	AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_163_), .C(rst_bF_buf59), .Y(_121__11_) );
	NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_12_), .B(_1004__bF_buf0), .Y(_168_) );
	AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_28_), .C(_1009__bF_buf2), .Y(_169_) );
	OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_146_), .C(_169_), .Y(_170_) );
	AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(biu_ahb_data_out_20_), .Y(_171_) );
	OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_171_), .C(_170_), .Y(_172_) );
	AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_168_), .C(rst_bF_buf58), .Y(_121__12_) );
	NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_13_), .B(_1004__bF_buf5), .Y(_173_) );
	AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_29_), .C(_1009__bF_buf1), .Y(_174_) );
	OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_146_), .C(_174_), .Y(_175_) );
	AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf1), .B(biu_ahb_data_out_21_), .Y(_176_) );
	OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_176_), .C(_175_), .Y(_177_) );
	AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_173_), .C(rst_bF_buf57), .Y(_121__13_) );
	NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_14_), .B(_1004__bF_buf4), .Y(_178_) );
	AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_30_), .C(_1009__bF_buf0), .Y(_179_) );
	OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_146_), .C(_179_), .Y(_180_) );
	NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_1004__bF_buf3), .Y(_181_) );
	OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_181_), .C(_180_), .Y(_182_) );
	AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_178_), .C(rst_bF_buf56), .Y(_121__14_) );
	NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .B(_1004__bF_buf2), .Y(_183_) );
	AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(biu_ahb_data_out_31_), .C(_1009__bF_buf3), .Y(_184_) );
	OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_146_), .C(_184_), .Y(_185_) );
	NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_1004__bF_buf1), .Y(_186_) );
	OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_186_), .C(_185_), .Y(_187_) );
	AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_183_), .C(rst_bF_buf55), .Y(_121__15_) );
	NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_16_), .B(_1004__bF_buf0), .Y(_188_) );
	OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_855_), .C(_1014_), .Y(_189_) );
	OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_116__1_), .B(_116__0_), .C(_189_), .Y(_190_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_16_), .B(_1031__bF_buf0), .C(_190_), .Y(_191_) );
	AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_188_), .C(rst_bF_buf54), .Y(_121__16_) );
	NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_17_), .B(_1004__bF_buf5), .Y(_192_) );
	NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_190_), .Y(_193_) );
	AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_192_), .C(rst_bF_buf53), .Y(_121__17_) );
	NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_18_), .B(_1004__bF_buf4), .Y(_194_) );
	NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_190_), .Y(_195_) );
	AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_194_), .C(rst_bF_buf52), .Y(_121__18_) );
	NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_19_), .B(_1004__bF_buf3), .Y(_196_) );
	NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_190_), .Y(_197_) );
	AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_196_), .C(rst_bF_buf51), .Y(_121__19_) );
	NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_20_), .B(_1004__bF_buf2), .Y(_198_) );
	NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_190_), .Y(_199_) );
	AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_198_), .C(rst_bF_buf50), .Y(_121__20_) );
	NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_21_), .B(_1004__bF_buf1), .Y(_200_) );
	NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_190_), .Y(_201_) );
	AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_200_), .C(rst_bF_buf49), .Y(_121__21_) );
	NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_22_), .B(_1004__bF_buf0), .Y(_202_) );
	NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_190_), .Y(_203_) );
	AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_202_), .C(rst_bF_buf48), .Y(_121__22_) );
	NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_23_), .B(_1004__bF_buf5), .Y(_204_) );
	NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_190_), .Y(_205_) );
	AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_204_), .C(rst_bF_buf47), .Y(_121__23_) );
	NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_24_), .B(_1004__bF_buf4), .Y(_206_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_24_), .B(_1031__bF_buf3), .C(_190_), .Y(_207_) );
	AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_206_), .C(rst_bF_buf46), .Y(_121__24_) );
	NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_25_), .B(_1004__bF_buf3), .Y(_208_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_25_), .B(_1031__bF_buf2), .C(_190_), .Y(_209_) );
	AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_208_), .C(rst_bF_buf45), .Y(_121__25_) );
	NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_26_), .B(_1004__bF_buf2), .Y(_210_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_26_), .B(_1031__bF_buf1), .C(_190_), .Y(_211_) );
	AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_210_), .C(rst_bF_buf44), .Y(_121__26_) );
	NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_27_), .B(_1004__bF_buf1), .Y(_212_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_27_), .B(_1031__bF_buf0), .C(_190_), .Y(_213_) );
	AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_212_), .C(rst_bF_buf43), .Y(_121__27_) );
	NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_28_), .B(_1004__bF_buf0), .Y(_214_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_28_), .B(_1031__bF_buf3), .C(_190_), .Y(_215_) );
	AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_214_), .C(rst_bF_buf42), .Y(_121__28_) );
	NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_29_), .B(_1004__bF_buf5), .Y(_216_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_29_), .B(_1031__bF_buf2), .C(_190_), .Y(_217_) );
	AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_216_), .C(rst_bF_buf41), .Y(_121__29_) );
	NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_30_), .B(_1004__bF_buf4), .Y(_218_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_30_), .B(_1031__bF_buf1), .C(_190_), .Y(_219_) );
	AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_218_), .C(rst_bF_buf40), .Y(_121__30_) );
	NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_31_), .B(_1004__bF_buf3), .Y(_220_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_31_), .B(_1031__bF_buf0), .C(_190_), .Y(_221_) );
	AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_220_), .C(rst_bF_buf39), .Y(_121__31_) );
	INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_0_), .Y(_222_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .C(biu_rdy_biu), .Y(_223_) );
	INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf38), .Y(_224_) );
	OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_0_), .B(_223__bF_buf7), .C(_224__bF_buf4), .Y(_225_) );
	AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223__bF_buf6), .C(_225_), .Y(_122__0_) );
	INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_1_), .Y(_226_) );
	OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_1_), .B(_223__bF_buf5), .C(_224__bF_buf3), .Y(_227_) );
	AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_223__bF_buf4), .C(_227_), .Y(_122__1_) );
	INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .Y(_228_) );
	OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_2_), .B(_223__bF_buf3), .C(_224__bF_buf2), .Y(_229_) );
	AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_223__bF_buf2), .C(_229_), .Y(_122__2_) );
	INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_3_), .Y(_230_) );
	OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_3_), .B(_223__bF_buf1), .C(_224__bF_buf1), .Y(_231_) );
	AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_223__bF_buf0), .C(_231_), .Y(_122__3_) );
	INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .Y(_232_) );
	OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_4_), .B(_223__bF_buf7), .C(_224__bF_buf0), .Y(_233_) );
	AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_223__bF_buf6), .C(_233_), .Y(_122__4_) );
	INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_5_), .Y(_234_) );
	OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_5_), .B(_223__bF_buf5), .C(_224__bF_buf4), .Y(_235_) );
	AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_223__bF_buf4), .C(_235_), .Y(_122__5_) );
	INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .Y(_236_) );
	OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_6_), .B(_223__bF_buf3), .C(_224__bF_buf3), .Y(_237_) );
	AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_223__bF_buf2), .C(_237_), .Y(_122__6_) );
	INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_7_), .Y(_238_) );
	OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_7_), .B(_223__bF_buf1), .C(_224__bF_buf2), .Y(_239_) );
	AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_223__bF_buf0), .C(_239_), .Y(_122__7_) );
	INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .Y(_240_) );
	OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_8_), .B(_223__bF_buf7), .C(_224__bF_buf1), .Y(_241_) );
	AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_223__bF_buf6), .C(_241_), .Y(_122__8_) );
	INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_9_), .Y(_242_) );
	OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_9_), .B(_223__bF_buf5), .C(_224__bF_buf0), .Y(_243_) );
	AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_223__bF_buf4), .C(_243_), .Y(_122__9_) );
	INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_10_), .Y(_244_) );
	OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_10_), .B(_223__bF_buf3), .C(_224__bF_buf4), .Y(_245_) );
	AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_223__bF_buf2), .C(_245_), .Y(_122__10_) );
	INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .Y(_246_) );
	OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_11_), .B(_223__bF_buf1), .C(_224__bF_buf3), .Y(_247_) );
	AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_223__bF_buf0), .C(_247_), .Y(_122__11_) );
	INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_12_), .Y(_248_) );
	OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_12_), .B(_223__bF_buf7), .C(_224__bF_buf2), .Y(_249_) );
	AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_223__bF_buf6), .C(_249_), .Y(_122__12_) );
	INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .Y(_250_) );
	OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_13_), .B(_223__bF_buf5), .C(_224__bF_buf1), .Y(_251_) );
	AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_223__bF_buf4), .C(_251_), .Y(_122__13_) );
	INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .Y(_252_) );
	OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_14_), .B(_223__bF_buf3), .C(_224__bF_buf0), .Y(_253_) );
	AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_223__bF_buf2), .C(_253_), .Y(_122__14_) );
	INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf6), .Y(_254_) );
	OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_15_), .B(_223__bF_buf1), .C(_224__bF_buf4), .Y(_255_) );
	AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_223__bF_buf0), .C(_255_), .Y(_122__15_) );
	INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_16_), .Y(_256_) );
	OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_16_), .B(_223__bF_buf7), .C(_224__bF_buf3), .Y(_257_) );
	AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_223__bF_buf6), .C(_257_), .Y(_122__16_) );
	INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_17_), .Y(_258_) );
	OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_17_), .B(_223__bF_buf5), .C(_224__bF_buf2), .Y(_259_) );
	AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_223__bF_buf4), .C(_259_), .Y(_122__17_) );
	INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .Y(_260_) );
	OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_18_), .B(_223__bF_buf3), .C(_224__bF_buf1), .Y(_261_) );
	AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_223__bF_buf2), .C(_261_), .Y(_122__18_) );
	INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_19_), .Y(_262_) );
	OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_19_), .B(_223__bF_buf1), .C(_224__bF_buf0), .Y(_263_) );
	AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_223__bF_buf0), .C(_263_), .Y(_122__19_) );
	INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf6), .Y(_264_) );
	OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_20_), .B(_223__bF_buf7), .C(_224__bF_buf4), .Y(_265_) );
	AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_223__bF_buf6), .C(_265_), .Y(_122__20_) );
	INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf3), .Y(_266_) );
	OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_21_), .B(_223__bF_buf5), .C(_224__bF_buf3), .Y(_267_) );
	AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_223__bF_buf4), .C(_267_), .Y(_122__21_) );
	INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf3), .Y(_268_) );
	OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_22_), .B(_223__bF_buf3), .C(_224__bF_buf2), .Y(_269_) );
	AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_223__bF_buf2), .C(_269_), .Y(_122__22_) );
	INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .Y(_270_) );
	OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_23_), .B(_223__bF_buf1), .C(_224__bF_buf1), .Y(_271_) );
	AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_223__bF_buf0), .C(_271_), .Y(_122__23_) );
	INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_272_) );
	OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_24_), .B(_223__bF_buf7), .C(_224__bF_buf0), .Y(_273_) );
	AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_223__bF_buf6), .C(_273_), .Y(_122__24_) );
	INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf3), .Y(_274_) );
	OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_25_), .B(_223__bF_buf5), .C(_224__bF_buf4), .Y(_275_) );
	AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_223__bF_buf4), .C(_275_), .Y(_122__25_) );
	INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf3), .Y(_276_) );
	OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_26_), .B(_223__bF_buf3), .C(_224__bF_buf3), .Y(_277_) );
	AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_223__bF_buf2), .C(_277_), .Y(_122__26_) );
	INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf3), .Y(_278_) );
	OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_27_), .B(_223__bF_buf1), .C(_224__bF_buf2), .Y(_279_) );
	AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_223__bF_buf0), .C(_279_), .Y(_122__27_) );
	INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf3), .Y(_280_) );
	OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_28_), .B(_223__bF_buf7), .C(_224__bF_buf1), .Y(_281_) );
	AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_223__bF_buf6), .C(_281_), .Y(_122__28_) );
	INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf3), .Y(_282_) );
	OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_29_), .B(_223__bF_buf5), .C(_224__bF_buf0), .Y(_283_) );
	AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_223__bF_buf4), .C(_283_), .Y(_122__29_) );
	INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf3), .Y(_284_) );
	OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_30_), .B(_223__bF_buf3), .C(_224__bF_buf4), .Y(_285_) );
	AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_223__bF_buf2), .C(_285_), .Y(_122__30_) );
	INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .Y(_286_) );
	OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_31_), .B(_223__bF_buf1), .C(_224__bF_buf3), .Y(_287_) );
	AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_223__bF_buf0), .C(_287_), .Y(_122__31_) );
	NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_698_), .Y(_288_) );
	INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_683_), .Y(_289_) );
	OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(addr_csr_0_), .C(_685_), .Y(_290_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(biu_exce_chk_opc_1_), .C(_688_), .Y(_291_) );
	AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_291_), .C(_693_), .Y(_292_) );
	NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_ahb_acc_fault), .B(gnd), .Y(_293_) );
	INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_293_), .Y(_294_) );
	NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_294_), .C(_292_), .Y(_295_) );
	OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(biu_ahb_rdy_ahb_bF_buf5), .C(_295_), .Y(_296_) );
	INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(_296_), .Y(_297_) );
	OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf1), .B(_288_), .C(_297_), .Y(_298_) );
	NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_698_), .Y(_299_) );
	NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_page_not_value), .B(_294_), .C(biu_addr_mis), .Y(_300_) );
	NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb_bF_buf4), .B(_629_), .Y(_301_) );
	NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_300_), .Y(_302_) );
	NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_698_), .Y(_303_) );
	NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(biu_rdy_biu), .B(_303_), .Y(_304_) );
	NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_955_), .Y(_305_) );
	INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_305_), .Y(_306_) );
	INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(_843_), .Y(_307_) );
	NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_695_), .Y(_308_) );
	INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_308_), .Y(_309_) );
	INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_649_), .Y(_310_) );
	NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_310_), .Y(_311_) );
	NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_310_), .Y(_312_) );
	INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_312_), .Y(_313_) );
	INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_954_), .Y(_314_) );
	NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_695_), .Y(_315_) );
	INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_315_), .Y(_316_) );
	NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_633_), .Y(_317_) );
	NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_956_), .Y(_318_) );
	OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_703_), .C(_654_), .Y(_319_) );
	OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_319_), .C(_297_), .Y(_320_) );
	NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_696_), .Y(_321_) );
	NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_705_), .Y(_322_) );
	NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_703_), .Y(_323_) );
	INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_323_), .Y(_324_) );
	OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_296_), .C(_629_), .Y(_325_) );
	AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_322_), .C(_321_), .D(_325_), .Y(_326_) );
	OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_326_), .C(_320_), .Y(_327_) );
	NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_705_), .Y(_328_) );
	INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_328_), .Y(_329_) );
	INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_330_) );
	NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_330_), .Y(_331_) );
	OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_329_), .C(_331_), .Y(_332_) );
	AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_316_), .C(_332_), .Y(_333_) );
	AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_302_), .C(_333_), .Y(_334_) );
	NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_652_), .Y(_335_) );
	INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_335_), .Y(_336_) );
	OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_702_), .C(_649_), .Y(_337_) );
	AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .C(_296_), .Y(_338_) );
	OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_334_), .C(_313_), .Y(_339_) );
	NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_310_), .Y(_340_) );
	NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_302_), .Y(_341_) );
	AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_340_), .C(_341_), .Y(_342_) );
	AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_342_), .C(_311_), .Y(_343_) );
	INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_311_), .Y(_344_) );
	NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_310_), .Y(_345_) );
	INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_844_), .Y(_346_) );
	OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_698_), .C(_346_), .Y(_347_) );
	OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_347_), .C(_297_), .Y(_348_) );
	OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_302_), .C(_348_), .Y(_349_) );
	OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_343_), .C(_309_), .Y(_350_) );
	NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_705_), .Y(_351_) );
	NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_302_), .Y(_352_) );
	AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_351_), .C(_352_), .Y(_353_) );
	AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_307_), .C(_353_), .D(_350_), .Y(_354_) );
	NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_694_), .Y(_355_) );
	NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_843_), .Y(_356_) );
	INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_356_), .Y(_357_) );
	OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_840_), .C(_357_), .Y(_358_) );
	OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_358_), .C(_297_), .Y(_359_) );
	OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_302_), .C(_359_), .Y(_360_) );
	NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_840_), .Y(_361_) );
	INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_362_) );
	OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_354_), .C(_362_), .Y(_363_) );
	NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_840_), .Y(_364_) );
	NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_302_), .Y(_365_) );
	AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_364_), .C(_365_), .Y(_366_) );
	AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_663_), .C(_366_), .D(_363_), .Y(_367_) );
	NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_694_), .Y(_368_) );
	NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_840_), .Y(_369_) );
	INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_369_), .Y(_370_) );
	OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_703_), .C(_370_), .Y(_371_) );
	OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_371_), .C(_297_), .Y(_372_) );
	OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_302_), .C(_372_), .Y(_373_) );
	OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_367_), .C(_306_), .Y(_374_) );
	NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_955_), .Y(_375_) );
	NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_302_), .Y(_376_) );
	AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_375_), .C(_376_), .Y(_377_) );
	AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_658_), .C(_377_), .D(_374_), .Y(_378_) );
	NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_955_), .Y(_379_) );
	INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_379_), .Y(_380_) );
	NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_955_), .Y(_381_) );
	OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_381_), .C(_297_), .Y(_382_) );
	OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_302_), .C(_382_), .Y(_383_) );
	OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_378_), .C(_304_), .Y(_384_) );
	NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_297_), .Y(_385_) );
	AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_302_), .C(_385_), .D(_384_), .Y(_386_) );
	NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_698_), .Y(_387_) );
	AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_387_), .C(_700_), .Y(_388_) );
	OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_386_), .C(_388_), .Y(_389_) );
	OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_297_), .C(_224__bF_buf2), .Y(_390_) );
	AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_298_), .C(_390_), .Y(_123__0_) );
	INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_387_), .Y(_391_) );
	INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_376_), .Y(_392_) );
	INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_365_), .Y(_393_) );
	INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_352_), .Y(_394_) );
	INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_341_), .Y(_395_) );
	NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_322_), .Y(_396_) );
	OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_330_), .C(_396_), .Y(_397_) );
	INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb_bF_buf3), .Y(_398_) );
	OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_mmu_st_page_fault), .B(biu_exce_chk_mmu_ld_page_fault), .C(biu_ahb_rdy_ahb_bF_buf2), .Y(_399_) );
	NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_300_), .Y(_400_) );
	AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_398_), .C(_400_), .Y(_401_) );
	NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(biu_exce_chk_opc_1_), .Y(_402_) );
	AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_673_), .C(_402_), .Y(_403_) );
	NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(addr_csr_0_), .Y(_404_) );
	NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(_686_), .C(_404_), .Y(_405_) );
	NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(biu_exce_chk_statu_cpu_2_), .C(_691_), .Y(_406_) );
	OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_406_), .Y(_407_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_293_), .C(_407_), .Y(_408_) );
	AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_398_), .C(_408_), .Y(_409_) );
	AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_409_), .C(_317_), .D(_401_), .Y(_410_) );
	OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_330_), .C(_329_), .Y(_411_) );
	AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_397_), .C(_411_), .Y(_412_) );
	INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_401_), .Y(_413_) );
	NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_409_), .Y(_414_) );
	OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_413_), .C(_414_), .Y(_415_) );
	OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_412_), .C(_313_), .Y(_416_) );
	AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_395_), .C(_340_), .Y(_417_) );
	NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_409_), .Y(_418_) );
	OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_413_), .C(_418_), .Y(_419_) );
	OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_417_), .C(_309_), .Y(_420_) );
	AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_394_), .C(_351_), .Y(_421_) );
	NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_409_), .Y(_422_) );
	OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_413_), .C(_422_), .Y(_423_) );
	OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_421_), .C(_362_), .Y(_424_) );
	AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_393_), .C(_364_), .Y(_425_) );
	NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_409_), .Y(_426_) );
	OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_413_), .C(_426_), .Y(_427_) );
	OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_425_), .C(_306_), .Y(_428_) );
	AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_392_), .C(_375_), .Y(_429_) );
	NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_409_), .Y(_430_) );
	OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_413_), .C(_430_), .Y(_431_) );
	OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf0), .B(biu_ahb_rdy_ahb_bF_buf1), .C(_295_), .Y(_432_) );
	AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_432_), .C(_299_), .D(_302_), .Y(_433_) );
	OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_429_), .C(_433_), .Y(_434_) );
	OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_401_), .C(_224__bF_buf1), .Y(_435_) );
	AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_391_), .C(_435_), .Y(_123__1_) );
	NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_955_), .Y(_436_) );
	INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_848_), .Y(_437_) );
	OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_703_), .C(biu_exce_chk_statu_biu_2_), .Y(_438_) );
	NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_703_), .Y(_439_) );
	INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_439_), .Y(_440_) );
	NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_310_), .Y(_441_) );
	INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_441_), .Y(_442_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_324_), .C(_442_), .Y(_443_) );
	NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_443_), .Y(_444_) );
	INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_445_) );
	OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(biu_ahb_rdy_ahb_bF_buf0), .C(_445_), .Y(_446_) );
	OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_695_), .C(_321_), .Y(_447_) );
	NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_447_), .Y(_448_) );
	AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_448_), .C(_446_), .Y(_449_) );
	OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_449_), .C(_437_), .Y(_450_) );
	INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_446_), .Y(_451_) );
	NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(_398_), .Y(_452_) );
	NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_408_), .Y(_453_) );
	AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_361_), .C(_453_), .Y(_454_) );
	AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_454_), .C(_436_), .Y(_455_) );
	NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_453_), .Y(_456_) );
	OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_446_), .C(_456_), .Y(_457_) );
	OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_455_), .C(_304_), .Y(_458_) );
	NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_453_), .Y(_459_) );
	NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_458_), .Y(_460_) );
	NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_446_), .Y(_461_) );
	OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_460_), .C(_461_), .Y(_462_) );
	NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf37), .B(_462_), .Y(_123__2_) );
	INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_31_), .Y(_463_) );
	INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mis), .Y(_464_) );
	INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .Y(_465_) );
	NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_693_), .Y(_466_) );
	INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_466_), .Y(_467_) );
	NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_467_), .Y(_468_) );
	NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_1014_), .Y(_469_) );
	INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_469_), .Y(_470_) );
	NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(biu_addr_mis), .Y(_471_) );
	INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_471_), .Y(_472_) );
	OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_472_), .C(_470_), .Y(_473_) );
	AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .C(_473_), .Y(_474_) );
	NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .Y(_475_) );
	NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .B(_693_), .Y(_476_) );
	NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_476_), .Y(_477_) );
	OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(biu_addr_mis), .C(_477_), .Y(_478_) );
	NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_687_), .Y(_479_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .C(_464_), .Y(_480_) );
	OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_472_), .C(_480_), .Y(_481_) );
	NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_481_), .Y(_482_) );
	AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_474_), .Y(_483_) );
	NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_638_), .Y(_484_) );
	INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_484_), .Y(_485_) );
	AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_641_), .C(_485_), .Y(_486_) );
	OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_483_), .C(_486_), .Y(_487_) );
	NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .B(_398_), .Y(_488_) );
	NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_408_), .Y(_489_) );
	NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_645__bF_buf0), .B(_661_), .Y(_490_) );
	OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf0), .B(_846_), .C(biu_exce_chk_statu_biu_3_), .Y(_491_) );
	NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_841_), .Y(_492_) );
	AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_492_), .C(_489_), .Y(_493_) );
	AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_493_), .C(rst_bF_buf36), .Y(_123__3_) );
	NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_432_), .Y(_494_) );
	OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf3), .B(biu_ahb_rdy_ahb_bF_buf5), .C(_445_), .Y(_495_) );
	INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_495_), .Y(_496_) );
	NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf2), .B(_398_), .Y(_497_) );
	OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_408_), .C(_702_), .Y(_498_) );
	OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_837__bF_buf3), .B(_496_), .C(_498_), .Y(_499_) );
	OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_842_), .C(_499_), .Y(_500_) );
	INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(_432_), .Y(_501_) );
	OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_658_), .C(_704_), .Y(_502_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_502_), .Y(_503_) );
	AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_654_), .C(_489_), .Y(_504_) );
	NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf1), .B(_304_), .Y(_505_) );
	NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_505_), .Y(_506_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_506_), .C(_500_), .Y(_507_) );
	AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_495_), .C(_459_), .D(_507_), .Y(_508_) );
	AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_387_), .C(_288_), .Y(_509_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_509_), .C(_508_), .Y(_510_) );
	INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_478_), .Y(_511_) );
	NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_472_), .Y(_512_) );
	INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_512_), .Y(_513_) );
	NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_513_), .Y(_514_) );
	NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_472_), .Y(_515_) );
	NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_31_), .B(_515_), .Y(_516_) );
	NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .Y(_517_) );
	MUX2X1 MUX2X1_58 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf0), .B(_463_), .S(_517_), .Y(_518_) );
	OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_518_), .C(_516_), .Y(_519_) );
	OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_1014_), .C(_519_), .Y(_520_) );
	OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_31_), .B(_470_), .C(_520_), .Y(_521_) );
	OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_480_), .C(_513_), .Y(_522_) );
	AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_480_), .C(_522_), .Y(_523_) );
	OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_523_), .C(_511_), .Y(_524_) );
	AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_463_), .C(_485_), .Y(_525_) );
	AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_501_), .C(_525_), .D(_524_), .Y(_526_) );
	AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_510_), .C(rst_bF_buf35), .Y(_123__4_) );
	INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_364_), .Y(_527_) );
	NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_453_), .Y(_528_) );
	INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_351_), .Y(_529_) );
	NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_453_), .Y(_530_) );
	NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_453_), .Y(_531_) );
	NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb_bF_buf4), .B(_635_), .Y(_532_) );
	AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(_654_), .C(_532_), .D(_295_), .Y(_533_) );
	OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_533_), .C(_531_), .Y(_534_) );
	INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_page_not_value), .Y(_535_) );
	OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_ahb_rdy_ahb_bF_buf3), .C(_399_), .Y(_536_) );
	INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_537_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_537_), .C(_295_), .Y(_538_) );
	AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_315_), .C(_328_), .Y(_539_) );
	AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_409_), .C(_539_), .D(_534_), .Y(_540_) );
	INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_538_), .Y(_541_) );
	OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_541_), .C(_336_), .Y(_542_) );
	AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_398_), .C(_408_), .Y(_543_) );
	INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_543_), .Y(_544_) );
	OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_544_), .C(_542_), .D(_540_), .Y(_545_) );
	INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_546_) );
	NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_295_), .Y(_547_) );
	AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_546_), .C(_441_), .Y(_548_) );
	AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_453_), .C(_548_), .D(_545_), .Y(_549_) );
	INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_550_) );
	OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_541_), .C(_550_), .Y(_551_) );
	OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_549_), .C(_418_), .Y(_552_) );
	INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_300_), .Y(_553_) );
	OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_553_), .C(_311_), .Y(_554_) );
	AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_345_), .C(_844_), .Y(_555_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_555_), .C(_552_), .Y(_556_) );
	AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_307_), .C(_530_), .D(_556_), .Y(_557_) );
	NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_538_), .Y(_558_) );
	OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_557_), .C(_529_), .Y(_559_) );
	AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_307_), .C(_422_), .D(_559_), .Y(_560_) );
	NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_538_), .Y(_561_) );
	OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_560_), .C(_357_), .Y(_562_) );
	NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_543_), .Y(_563_) );
	AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_663_), .C(_563_), .D(_562_), .Y(_564_) );
	INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_841_), .Y(_565_) );
	NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_565_), .Y(_566_) );
	OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_564_), .C(_437_), .Y(_567_) );
	AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_696_), .C(_528_), .D(_567_), .Y(_568_) );
	NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_538_), .Y(_569_) );
	OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_568_), .C(_527_), .Y(_570_) );
	AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_663_), .C(_426_), .D(_570_), .Y(_571_) );
	NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_538_), .Y(_572_) );
	OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_571_), .C(_370_), .Y(_573_) );
	OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(biu_addr_mis), .C(_484_), .Y(_574_) );
	INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_574_), .Y(_575_) );
	INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_514_), .Y(_576_) );
	NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(_517_), .Y(_577_) );
	OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_517_), .C(_577_), .Y(_578_) );
	AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_31_), .B(_469_), .C(_481_), .Y(_579_) );
	OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_578_), .C(_579_), .Y(_580_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_580_), .C(_576_), .Y(_581_) );
	NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_544_), .Y(_582_) );
	AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_575_), .C(_582_), .Y(_583_) );
	AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_583_), .C(rst_bF_buf34), .Y(_123__5_) );
	OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf3), .B(biu_ahb_rdy_ahb_bF_buf2), .C(_399_), .Y(_584_) );
	OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_553_), .C(_379_), .Y(_585_) );
	INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_582_), .Y(_586_) );
	NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_409_), .Y(_587_) );
	INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_584_), .Y(_588_) );
	AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_588_), .C(_321_), .Y(_589_) );
	INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_322_), .Y(_590_) );
	OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_408_), .C(_323_), .Y(_591_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf2), .B(_590_), .C(_591_), .Y(_592_) );
	OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_589_), .C(_587_), .Y(_593_) );
	OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_553_), .C(_317_), .Y(_594_) );
	OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf1), .B(biu_ahb_rdy_ahb_bF_buf1), .C(_295_), .Y(_595_) );
	AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_318_), .C(_844_), .Y(_596_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_596_), .C(_593_), .Y(_597_) );
	AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_307_), .C(_530_), .D(_597_), .Y(_598_) );
	OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_598_), .C(_529_), .Y(_599_) );
	AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_307_), .C(_422_), .D(_599_), .Y(_600_) );
	OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_600_), .C(_357_), .Y(_601_) );
	AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_663_), .C(_563_), .D(_601_), .Y(_602_) );
	OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_602_), .C(_437_), .Y(_603_) );
	AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_696_), .C(_528_), .D(_603_), .Y(_604_) );
	OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_604_), .C(_527_), .Y(_605_) );
	AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_663_), .C(_426_), .D(_605_), .Y(_606_) );
	OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_606_), .C(_370_), .Y(_607_) );
	NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_607_), .Y(_608_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf0), .B(_398_), .C(_295_), .Y(_609_) );
	AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_847_), .C(_436_), .Y(_610_) );
	AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_453_), .C(_610_), .D(_608_), .Y(_611_) );
	INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_375_), .Y(_612_) );
	OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_496_), .C(_612_), .Y(_613_) );
	OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_611_), .C(_430_), .Y(_614_) );
	AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_381_), .C(_957_), .Y(_615_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_615_), .C(_614_), .Y(_616_) );
	NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf3), .B(_474_), .Y(_617_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_579_), .C(_617_), .Y(_618_) );
	NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_609_), .Y(_619_) );
	AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_575_), .C(_619_), .Y(_620_) );
	AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_620_), .C(rst_bF_buf33), .Y(_123__6_) );
	NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_464_), .Y(_621_) );
	NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_621_), .Y(_622_) );
	INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_622_), .Y(_623_) );
	NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_961_), .Y(_624_) );
	NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_624_), .Y(biu_ahb_w32) );
	NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_623_), .Y(biu_ahb_w16) );
	NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_623_), .Y(biu_ahb_w8) );
	NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_635_), .Y(_625_) );
	OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_698_), .C(_442_), .Y(_626_) );
	AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_625_), .C(_626_), .Y(_627_) );
	AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_627_), .C(_623_), .Y(biu_ahb_r32) );
	AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_440_), .C(_623_), .Y(biu_ahb_r16) );
	AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_324_), .C(_623_), .Y(biu_ahb_r8) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_121__0_), .Q(biu_biu_data_out_0_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_121__1_), .Q(biu_biu_data_out_1_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_121__2_), .Q(biu_biu_data_out_2_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_121__3_), .Q(biu_biu_data_out_3_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_121__4_), .Q(biu_biu_data_out_4_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_121__5_), .Q(biu_biu_data_out_5_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_121__6_), .Q(biu_biu_data_out_6_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_121__7_), .Q(biu_biu_data_out_7_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_121__8_), .Q(biu_biu_data_out_8_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_121__9_), .Q(biu_biu_data_out_9_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_121__10_), .Q(biu_biu_data_out_10_) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_121__11_), .Q(biu_biu_data_out_11_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_121__12_), .Q(biu_biu_data_out_12_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_121__13_), .Q(biu_biu_data_out_13_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_121__14_), .Q(biu_biu_data_out_14_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_121__15_), .Q(biu_biu_data_out_15_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_121__16_), .Q(biu_biu_data_out_16_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_121__17_), .Q(biu_biu_data_out_17_) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_121__18_), .Q(biu_biu_data_out_18_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_121__19_), .Q(biu_biu_data_out_19_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_121__20_), .Q(biu_biu_data_out_20_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_121__21_), .Q(biu_biu_data_out_21_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_121__22_), .Q(biu_biu_data_out_22_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_121__23_), .Q(biu_biu_data_out_23_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_121__24_), .Q(biu_biu_data_out_24_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_121__25_), .Q(biu_biu_data_out_25_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_121__26_), .Q(biu_biu_data_out_26_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_121__27_), .Q(biu_biu_data_out_27_) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_121__28_), .Q(biu_biu_data_out_28_) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_121__29_), .Q(biu_biu_data_out_29_) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_121__30_), .Q(biu_biu_data_out_30_) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_121__31_), .Q(biu_biu_data_out_31_) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_122__0_), .Q(biu_ins_0_) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_122__1_), .Q(biu_ins_1_) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_122__2_), .Q(biu_ins_2_) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_122__3_), .Q(biu_ins_3_) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_122__4_), .Q(biu_ins_4_) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_122__5_), .Q(biu_ins_5_) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_122__6_), .Q(biu_ins_6_) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_122__7_), .Q(biu_ins_7_) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_122__8_), .Q(biu_ins_8_) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_122__9_), .Q(biu_ins_9_) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_122__10_), .Q(biu_ins_10_) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_122__11_), .Q(biu_ins_11_) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_122__12_), .Q(biu_ins_12_) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_122__13_), .Q(biu_ins_13_) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_122__14_), .Q(biu_ins_14_) );
	DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_122__15_), .Q(biu_ins_15_) );
	DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_122__16_), .Q(biu_ins_16_) );
	DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_122__17_), .Q(biu_ins_17_) );
	DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_122__18_), .Q(biu_ins_18_) );
	DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_122__19_), .Q(biu_ins_19_) );
	DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_122__20_), .Q(biu_ins_20_) );
	DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_122__21_), .Q(biu_ins_21_) );
	DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_122__22_), .Q(biu_ins_22_) );
	DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_122__23_), .Q(biu_ins_23_) );
	DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_122__24_), .Q(biu_ins_24_) );
	DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_122__25_), .Q(biu_ins_25_) );
	DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_122__26_), .Q(biu_ins_26_) );
	DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_122__27_), .Q(biu_ins_27_) );
	DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_122__28_), .Q(biu_ins_28_) );
	DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_122__29_), .Q(biu_ins_29_) );
	DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_122__30_), .Q(biu_ins_30_) );
	DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_122__31_), .Q(biu_ins_31_) );
	DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_123__0_), .Q(biu_exce_chk_statu_biu_0_) );
	DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_123__1_), .Q(biu_exce_chk_statu_biu_1_) );
	DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_123__2_), .Q(biu_exce_chk_statu_biu_2_) );
	DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_123__3_), .Q(biu_exce_chk_statu_biu_3_) );
	DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_123__4_), .Q(biu_exce_chk_statu_biu_4_) );
	DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_123__5_), .Q(biu_exce_chk_statu_biu_5_) );
	DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_123__6_), .Q(biu_exce_chk_statu_biu_6_) );
	AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_in_0_), .B(biu_ahb_statu_ahb_bF_buf4), .Y(_119__0_) );
	AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_1_), .Y(_119__1_) );
	AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_2_), .Y(_119__2_) );
	AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_3_), .Y(_119__3_) );
	AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_4_), .Y(_119__4_) );
	AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_5_), .Y(_119__5_) );
	AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_6_), .Y(_119__6_) );
	AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_7_), .Y(_119__7_) );
	AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_8_), .Y(_119__8_) );
	AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_9_), .Y(_119__9_) );
	AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_10_), .Y(_119__10_) );
	AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_11_), .Y(_119__11_) );
	AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_12_), .Y(_119__12_) );
	AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_13_), .Y(_119__13_) );
	AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_14_), .Y(_119__14_) );
	AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_15_), .Y(_119__15_) );
	AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_16_), .Y(_119__16_) );
	AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_17_), .Y(_119__17_) );
	AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_18_), .Y(_119__18_) );
	AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_19_), .Y(_119__19_) );
	AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_20_), .Y(_119__20_) );
	AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_21_), .Y(_119__21_) );
	AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_22_), .Y(_119__22_) );
	AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_23_), .Y(_119__23_) );
	AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_24_), .Y(_119__24_) );
	AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_25_), .Y(_119__25_) );
	AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_26_), .Y(_119__26_) );
	AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .B(biu_ahb_data_in_27_), .Y(_119__27_) );
	AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(biu_ahb_data_in_28_), .Y(_119__28_) );
	AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf0), .B(biu_ahb_data_in_29_), .Y(_119__29_) );
	AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf4), .B(biu_ahb_data_in_30_), .Y(_119__30_) );
	AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf3), .B(biu_ahb_data_in_31_), .Y(_119__31_) );
	INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf2), .Y(_1067_) );
	INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(hready), .Y(_1068_) );
	NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf4), .Y(biu_ahb_rdy_ahb) );
	NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(hrdata[0]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1069_) );
	OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_0_), .Y(_1070_) );
	AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1070_), .C(rst_bF_buf32), .Y(_1065__0_) );
	NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(hrdata[1]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1071_) );
	OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_1_), .Y(_1072_) );
	AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1072_), .C(rst_bF_buf31), .Y(_1065__1_) );
	NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(hrdata[2]), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1073_) );
	OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_2_), .Y(_1074_) );
	AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1074_), .C(rst_bF_buf30), .Y(_1065__2_) );
	NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(hrdata[3]), .B(biu_ahb_rdy_ahb_bF_buf3), .Y(_1075_) );
	OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_3_), .Y(_1076_) );
	AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1076_), .C(rst_bF_buf29), .Y(_1065__3_) );
	NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(hrdata[4]), .B(biu_ahb_rdy_ahb_bF_buf2), .Y(_1077_) );
	OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_4_), .Y(_1078_) );
	AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1078_), .C(rst_bF_buf28), .Y(_1065__4_) );
	NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(hrdata[5]), .B(biu_ahb_rdy_ahb_bF_buf1), .Y(_1079_) );
	OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_5_), .Y(_1080_) );
	AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(_1080_), .C(rst_bF_buf27), .Y(_1065__5_) );
	NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(hrdata[6]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1081_) );
	OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_6_), .Y(_1082_) );
	AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1082_), .C(rst_bF_buf26), .Y(_1065__6_) );
	NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(hrdata[7]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1083_) );
	OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_7_), .Y(_1084_) );
	AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1084_), .C(rst_bF_buf25), .Y(_1065__7_) );
	NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(hrdata[8]), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1085_) );
	OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_8_), .Y(_1086_) );
	AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1086_), .C(rst_bF_buf24), .Y(_1065__8_) );
	NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(hrdata[9]), .B(biu_ahb_rdy_ahb_bF_buf3), .Y(_1087_) );
	OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_9_), .Y(_1088_) );
	AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(_1088_), .C(rst_bF_buf23), .Y(_1065__9_) );
	NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(hrdata[10]), .B(biu_ahb_rdy_ahb_bF_buf2), .Y(_1089_) );
	OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_10_), .Y(_1090_) );
	AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1090_), .C(rst_bF_buf22), .Y(_1065__10_) );
	NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(hrdata[11]), .B(biu_ahb_rdy_ahb_bF_buf1), .Y(_1091_) );
	OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_11_), .Y(_1092_) );
	AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(_1092_), .C(rst_bF_buf21), .Y(_1065__11_) );
	NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(hrdata[12]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1093_) );
	OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_12_), .Y(_1094_) );
	AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1094_), .C(rst_bF_buf20), .Y(_1065__12_) );
	NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(hrdata[13]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1095_) );
	OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_13_), .Y(_1096_) );
	AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1096_), .C(rst_bF_buf19), .Y(_1065__13_) );
	NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(hrdata[14]), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1097_) );
	OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_14_), .Y(_1098_) );
	AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1098_), .C(rst_bF_buf18), .Y(_1065__14_) );
	NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(hrdata[15]), .B(biu_ahb_rdy_ahb_bF_buf3), .Y(_1099_) );
	OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_15_), .Y(_1100_) );
	AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1100_), .C(rst_bF_buf17), .Y(_1065__15_) );
	NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(hrdata[16]), .B(biu_ahb_rdy_ahb_bF_buf2), .Y(_1101_) );
	OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_16_), .Y(_1102_) );
	AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(_1102_), .C(rst_bF_buf16), .Y(_1065__16_) );
	NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(hrdata[17]), .B(biu_ahb_rdy_ahb_bF_buf1), .Y(_1103_) );
	OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_17_), .Y(_1104_) );
	AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1104_), .C(rst_bF_buf15), .Y(_1065__17_) );
	NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(hrdata[18]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1105_) );
	OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_18_), .Y(_1106_) );
	AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1106_), .C(rst_bF_buf14), .Y(_1065__18_) );
	NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(hrdata[19]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1107_) );
	OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_19_), .Y(_1108_) );
	AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_1108_), .C(rst_bF_buf13), .Y(_1065__19_) );
	NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(hrdata[20]), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1109_) );
	OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_20_), .Y(_1110_) );
	AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1109_), .B(_1110_), .C(rst_bF_buf12), .Y(_1065__20_) );
	NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(hrdata[21]), .B(biu_ahb_rdy_ahb_bF_buf3), .Y(_1111_) );
	OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_21_), .Y(_1112_) );
	AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .B(_1112_), .C(rst_bF_buf11), .Y(_1065__21_) );
	NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(hrdata[22]), .B(biu_ahb_rdy_ahb_bF_buf2), .Y(_1113_) );
	OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_22_), .Y(_1114_) );
	AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .B(_1114_), .C(rst_bF_buf10), .Y(_1065__22_) );
	NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(hrdata[23]), .B(biu_ahb_rdy_ahb_bF_buf1), .Y(_1115_) );
	OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_23_), .Y(_1116_) );
	AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1116_), .C(rst_bF_buf9), .Y(_1065__23_) );
	NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(hrdata[24]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1117_) );
	OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_24_), .Y(_1118_) );
	AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1118_), .C(rst_bF_buf8), .Y(_1065__24_) );
	NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(hrdata[25]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1119_) );
	OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_25_), .Y(_1120_) );
	AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_1120_), .C(rst_bF_buf7), .Y(_1065__25_) );
	NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(hrdata[26]), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1121_) );
	OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_26_), .Y(_1122_) );
	AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1122_), .C(rst_bF_buf6), .Y(_1065__26_) );
	NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(hrdata[27]), .B(biu_ahb_rdy_ahb_bF_buf3), .Y(_1123_) );
	OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1068__bF_buf1), .C(biu_ahb_data_ahb_27_), .Y(_1124_) );
	AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .C(rst_bF_buf5), .Y(_1065__27_) );
	NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(hrdata[28]), .B(biu_ahb_rdy_ahb_bF_buf2), .Y(_1125_) );
	OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1068__bF_buf0), .C(biu_ahb_data_ahb_28_), .Y(_1126_) );
	AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(_1126_), .C(rst_bF_buf4), .Y(_1065__28_) );
	NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(hrdata[29]), .B(biu_ahb_rdy_ahb_bF_buf1), .Y(_1127_) );
	OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1068__bF_buf4), .C(biu_ahb_data_ahb_29_), .Y(_1128_) );
	AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1128_), .C(rst_bF_buf3), .Y(_1065__29_) );
	NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(hrdata[30]), .B(biu_ahb_rdy_ahb_bF_buf0), .Y(_1129_) );
	OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1068__bF_buf3), .C(biu_ahb_data_ahb_30_), .Y(_1130_) );
	AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1130_), .C(rst_bF_buf2), .Y(_1065__30_) );
	NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(hrdata[31]), .B(biu_ahb_rdy_ahb_bF_buf5), .Y(_1131_) );
	OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1068__bF_buf2), .C(biu_ahb_data_ahb_31_), .Y(_1132_) );
	AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1132_), .C(rst_bF_buf1), .Y(_1065__31_) );
	INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_w32), .Y(_1133_) );
	INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_w8), .Y(_1134_) );
	INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_w16), .Y(_1135_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1134_), .C(_1135_), .Y(_1136_) );
	INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_r16), .Y(_1137_) );
	INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_r32), .Y(_1138_) );
	INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_r8), .Y(_1139_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1138_), .C(_1139_), .Y(_1140_) );
	OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1140_), .C(_1067__bF_buf2), .Y(_1141_) );
	INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(hresp), .Y(_1142_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_statu_ahb_bF_buf1), .B(_1068__bF_buf1), .C(_1142_), .Y(_1143_) );
	AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1143_), .C(rst_bF_buf0), .Y(_1066_) );
	AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1067__bF_buf1), .Y(_120_) );
	NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1133_), .Y(_117__1_) );
	NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1135_), .Y(_117__0_) );
	INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_118__1_) );
	NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1142_), .Y(biu_ahb_ahb_acc_fault) );
	INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_0_), .Y(_1144_) );
	NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1069_), .Y(biu_ahb_data_out_0_) );
	INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_1_), .Y(_1145_) );
	NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_1071_), .Y(biu_ahb_data_out_1_) );
	INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_2_), .Y(_1146_) );
	NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_1073_), .Y(biu_ahb_data_out_2_) );
	INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_3_), .Y(_1147_) );
	NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1075_), .Y(biu_ahb_data_out_3_) );
	INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_4_), .Y(_1148_) );
	NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1077_), .Y(biu_ahb_data_out_4_) );
	INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_5_), .Y(_1149_) );
	NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_1079_), .Y(biu_ahb_data_out_5_) );
	INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_6_), .Y(_1150_) );
	NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1081_), .Y(biu_ahb_data_out_6_) );
	INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_7_), .Y(_1151_) );
	NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1083_), .Y(biu_ahb_data_out_7_) );
	INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_8_), .Y(_1152_) );
	NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_1085_), .Y(biu_ahb_data_out_8_) );
	INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_9_), .Y(_1153_) );
	NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1087_), .Y(biu_ahb_data_out_9_) );
	INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_10_), .Y(_1154_) );
	NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .B(_1089_), .Y(biu_ahb_data_out_10_) );
	INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_11_), .Y(_1155_) );
	NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1091_), .Y(biu_ahb_data_out_11_) );
	INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_12_), .Y(_1156_) );
	NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .B(_1093_), .Y(biu_ahb_data_out_12_) );
	INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_13_), .Y(_1157_) );
	NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1095_), .Y(biu_ahb_data_out_13_) );
	INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_14_), .Y(_1158_) );
	NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .B(_1097_), .Y(biu_ahb_data_out_14_) );
	INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_15_), .Y(_1159_) );
	NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1099_), .Y(biu_ahb_data_out_15_) );
	INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_16_), .Y(_1160_) );
	NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1101_), .Y(biu_ahb_data_out_16_) );
	INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_17_), .Y(_1161_) );
	NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(_1103_), .Y(biu_ahb_data_out_17_) );
	INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_18_), .Y(_1162_) );
	NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_1105_), .Y(biu_ahb_data_out_18_) );
	INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_19_), .Y(_1163_) );
	NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1107_), .Y(biu_ahb_data_out_19_) );
	INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_20_), .Y(_1164_) );
	NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1109_), .Y(biu_ahb_data_out_20_) );
	INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_21_), .Y(_1165_) );
	NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1111_), .Y(biu_ahb_data_out_21_) );
	INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_22_), .Y(_1166_) );
	NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1113_), .Y(biu_ahb_data_out_22_) );
	INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_23_), .Y(_1167_) );
	NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_1115_), .Y(biu_ahb_data_out_23_) );
	INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_24_), .Y(_1168_) );
	NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1117_), .Y(biu_ahb_data_out_24_) );
	INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_25_), .Y(_1169_) );
	NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1119_), .Y(biu_ahb_data_out_25_) );
	INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_26_), .Y(_1170_) );
	NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1121_), .Y(biu_ahb_data_out_26_) );
	INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_27_), .Y(_1171_) );
	NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1123_), .Y(biu_ahb_data_out_27_) );
	INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_28_), .Y(_1172_) );
	NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_1125_), .Y(biu_ahb_data_out_28_) );
	INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_29_), .Y(_1173_) );
	NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1127_), .Y(biu_ahb_data_out_29_) );
	INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_30_), .Y(_1174_) );
	NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_1129_), .Y(biu_ahb_data_out_30_) );
	INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_ahb_31_), .Y(_1175_) );
	NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1131_), .Y(biu_ahb_data_out_31_) );
	DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_1065__0_), .Q(biu_ahb_data_ahb_0_) );
	DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_1065__1_), .Q(biu_ahb_data_ahb_1_) );
	DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1065__2_), .Q(biu_ahb_data_ahb_2_) );
	DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_1065__3_), .Q(biu_ahb_data_ahb_3_) );
	DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1065__4_), .Q(biu_ahb_data_ahb_4_) );
	DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1065__5_), .Q(biu_ahb_data_ahb_5_) );
	DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1065__6_), .Q(biu_ahb_data_ahb_6_) );
	DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1065__7_), .Q(biu_ahb_data_ahb_7_) );
	DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1065__8_), .Q(biu_ahb_data_ahb_8_) );
	DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1065__9_), .Q(biu_ahb_data_ahb_9_) );
	DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1065__10_), .Q(biu_ahb_data_ahb_10_) );
	DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1065__11_), .Q(biu_ahb_data_ahb_11_) );
	DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1065__12_), .Q(biu_ahb_data_ahb_12_) );
	DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1065__13_), .Q(biu_ahb_data_ahb_13_) );
	DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1065__14_), .Q(biu_ahb_data_ahb_14_) );
	DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1065__15_), .Q(biu_ahb_data_ahb_15_) );
	DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1065__16_), .Q(biu_ahb_data_ahb_16_) );
	DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1065__17_), .Q(biu_ahb_data_ahb_17_) );
	DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1065__18_), .Q(biu_ahb_data_ahb_18_) );
	DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1065__19_), .Q(biu_ahb_data_ahb_19_) );
	DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1065__20_), .Q(biu_ahb_data_ahb_20_) );
	DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1065__21_), .Q(biu_ahb_data_ahb_21_) );
	DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1065__22_), .Q(biu_ahb_data_ahb_22_) );
	DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1065__23_), .Q(biu_ahb_data_ahb_23_) );
	DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1065__24_), .Q(biu_ahb_data_ahb_24_) );
	DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1065__25_), .Q(biu_ahb_data_ahb_25_) );
	DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1065__26_), .Q(biu_ahb_data_ahb_26_) );
	DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1065__27_), .Q(biu_ahb_data_ahb_27_) );
	DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1065__28_), .Q(biu_ahb_data_ahb_28_) );
	DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1065__29_), .Q(biu_ahb_data_ahb_29_) );
	DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1065__30_), .Q(biu_ahb_data_ahb_30_) );
	DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1065__31_), .Q(biu_ahb_data_ahb_31_) );
	DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1066_), .Q(biu_ahb_statu_ahb) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(biu_exce_chk_statu_cpu_0_), .Y(_1176_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_1_), .Y(_1177_) );
	NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1177_), .Y(_1178_) );
	NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mis), .B(_1178_), .Y(_1179_) );
	INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .Y(biu_exce_chk_ins_addr_mis) );
	INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1180_) );
	NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(biu_ahb_ahb_acc_fault), .Y(_1181_) );
	NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1180_), .Y(biu_exce_chk_ins_acc_fault) );
	INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .Y(_1182_) );
	INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .Y(_1183_) );
	NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1176_), .Y(_1184_) );
	NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mis), .B(_1184_), .Y(_1185_) );
	NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1185_), .Y(biu_exce_chk_load_addr_mis) );
	NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1181_), .C(_1176_), .Y(_1186_) );
	INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .Y(_1187_) );
	NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(biu_exce_chk_statu_biu_0_), .Y(_1188_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .B(_1187_), .C(_1188_), .Y(_1189_) );
	INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf2), .Y(_1190_) );
	INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .Y(_1191_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf3), .B(_1190_), .C(_1191_), .Y(_1192_) );
	INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .Y(_1193_) );
	NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(biu_exce_chk_statu_biu_2_), .C(_1188_), .Y(_1194_) );
	NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_exce_chk_statu_biu_4_bF_buf2), .Y(_1195_) );
	NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf1), .B(_1195_), .Y(_1196_) );
	OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1189_), .C(_1194_), .D(_1196_), .Y(_1197_) );
	NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1197_), .Y(_1198_) );
	NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf0), .B(_1191_), .Y(_1199_) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(biu_exce_chk_statu_biu_0_), .Y(_1200_) );
	NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .B(_1187_), .Y(_1201_) );
	NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(_1193_), .Y(_1202_) );
	AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1202_), .C(_1200_), .Y(_1203_) );
	NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_1203_), .C(_1186_), .Y(_1204_) );
	NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1198_), .Y(biu_exce_chk_load_acc_fault) );
	NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .B(_1185_), .Y(biu_exce_chk_st_addr_mis) );
	OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_exce_chk_statu_biu_4_bF_buf1), .C(biu_exce_chk_statu_biu_6_bF_buf3), .Y(_1205_) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1190_), .Y(_1206_) );
	AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_exce_chk_statu_biu_4_bF_buf0), .Y(_1207_) );
	NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_6_bF_buf2), .B(biu_exce_chk_statu_biu_5_), .C(biu_exce_chk_statu_biu_4_bF_buf3), .Y(_1208_) );
	OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1202_), .C(_1207_), .D(_1208_), .Y(_1209_) );
	NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_1186_), .C(_1209_), .Y(_1210_) );
	AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1206_), .C(_1210_), .Y(biu_exce_chk_st_acc_fault) );
	AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_mmu_ld_page_fault), .B(biu_ahb_rdy_ahb_bF_buf4), .Y(_1211_) );
	NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(_1193_), .Y(_1212_) );
	NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(_1212_), .Y(_1213_) );
	OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_page_not_value), .B(_1211_), .C(_1213_), .Y(_1214_) );
	NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1214_), .Y(biu_exce_chk_ins_page_fault) );
	INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .Y(_1215_) );
	AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_1215_), .C(_1214_), .Y(biu_exce_chk_ld_page_fault) );
	INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .Y(_1216_) );
	AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_rdy_ahb_bF_buf3), .B(biu_exce_chk_mmu_st_page_fault), .C(biu_exce_chk_page_not_value), .Y(_1217_) );
	NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1217_), .C(_1216_), .Y(biu_exce_chk_st_page_fault) );
	INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .Y(_1220_) );
	NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(biu_exce_chk_statu_biu_1_), .Y(_1221_) );
	INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(_1221__bF_buf4), .Y(_1222_) );
	OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag1_0_), .Y(_1223_) );
	AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1221__bF_buf3), .B(_1220__bF_buf4), .C(rst_bF_buf70), .Y(_1224_) );
	INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_1224__bF_buf3), .Y(_1225_) );
	NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1225__bF_buf5), .Y(_1218__0_) );
	OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag1_1_), .Y(_1226_) );
	NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1225__bF_buf4), .Y(_1218__1_) );
	INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_2_), .Y(_1227_) );
	NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(_1221__bF_buf2), .Y(_1228_) );
	OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_12_), .B(_1228__bF_buf5), .C(_1224__bF_buf2), .Y(_1229_) );
	AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .B(_1228__bF_buf4), .C(_1229_), .Y(_1218__2_) );
	INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_3_), .Y(_1230_) );
	OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_13_), .B(_1228__bF_buf3), .C(_1224__bF_buf1), .Y(_1231_) );
	AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1228__bF_buf2), .C(_1231_), .Y(_1218__3_) );
	INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_4_), .Y(_1232_) );
	OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_14_), .B(_1228__bF_buf1), .C(_1224__bF_buf0), .Y(_1233_) );
	AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1228__bF_buf0), .C(_1233_), .Y(_1218__4_) );
	INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_5_), .Y(_1234_) );
	OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_15_), .B(_1228__bF_buf5), .C(_1224__bF_buf3), .Y(_1235_) );
	AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1228__bF_buf4), .C(_1235_), .Y(_1218__5_) );
	INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_6_), .Y(_1236_) );
	OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_16_), .B(_1228__bF_buf3), .C(_1224__bF_buf2), .Y(_1237_) );
	AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1228__bF_buf2), .C(_1237_), .Y(_1218__6_) );
	INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_7_), .Y(_1238_) );
	OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_17_), .B(_1228__bF_buf1), .C(_1224__bF_buf1), .Y(_1239_) );
	AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1228__bF_buf0), .C(_1239_), .Y(_1218__7_) );
	INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_8_), .Y(_1240_) );
	OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_18_), .B(_1228__bF_buf5), .C(_1224__bF_buf0), .Y(_1241_) );
	AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_1228__bF_buf4), .C(_1241_), .Y(_1218__8_) );
	INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_9_), .Y(_1242_) );
	OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_19_), .B(_1228__bF_buf3), .C(_1224__bF_buf3), .Y(_1243_) );
	AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_1228__bF_buf2), .C(_1243_), .Y(_1218__9_) );
	INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_10_), .Y(_1244_) );
	OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_20_), .B(_1228__bF_buf1), .C(_1224__bF_buf2), .Y(_1245_) );
	AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1228__bF_buf0), .C(_1245_), .Y(_1218__10_) );
	INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_11_), .Y(_1246_) );
	OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_21_), .B(_1228__bF_buf5), .C(_1224__bF_buf1), .Y(_1247_) );
	AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1228__bF_buf4), .C(_1247_), .Y(_1218__11_) );
	OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag1_12_), .Y(_1248_) );
	INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(_1228__bF_buf3), .Y(_1249_) );
	NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_10_), .B(_1249__bF_buf3), .Y(_1250_) );
	AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1248_), .C(_1225__bF_buf3), .Y(_1218__12_) );
	OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag1_13_), .Y(_1251_) );
	NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_11_), .B(_1249__bF_buf2), .Y(_1252_) );
	AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1251_), .C(_1225__bF_buf2), .Y(_1218__13_) );
	OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag1_14_), .Y(_1253_) );
	NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_12_), .B(_1249__bF_buf1), .Y(_1254_) );
	AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1253_), .C(_1225__bF_buf1), .Y(_1218__14_) );
	OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag1_15_), .Y(_1255_) );
	NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_13_), .B(_1249__bF_buf0), .Y(_1256_) );
	AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1255_), .C(_1225__bF_buf0), .Y(_1218__15_) );
	OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag1_16_), .Y(_1257_) );
	NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_14_), .B(_1249__bF_buf3), .Y(_1258_) );
	AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_1257_), .C(_1225__bF_buf5), .Y(_1218__16_) );
	OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag1_17_), .Y(_1259_) );
	NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_15_), .B(_1249__bF_buf2), .Y(_1260_) );
	AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1259_), .C(_1225__bF_buf4), .Y(_1218__17_) );
	OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag1_18_), .Y(_1261_) );
	NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_16_), .B(_1249__bF_buf1), .Y(_1262_) );
	AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1261_), .C(_1225__bF_buf3), .Y(_1218__18_) );
	OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag1_19_), .Y(_1263_) );
	NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_17_), .B(_1249__bF_buf0), .Y(_1264_) );
	AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1263_), .C(_1225__bF_buf2), .Y(_1218__19_) );
	OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag1_20_), .Y(_1265_) );
	NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_18_), .B(_1249__bF_buf3), .Y(_1266_) );
	AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1265_), .C(_1225__bF_buf1), .Y(_1218__20_) );
	OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag1_21_), .Y(_1267_) );
	NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_19_), .B(_1249__bF_buf2), .Y(_1268_) );
	AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1267_), .C(_1225__bF_buf0), .Y(_1218__21_) );
	OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag1_22_), .Y(_1269_) );
	NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_20_), .B(_1249__bF_buf1), .Y(_1270_) );
	AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1269_), .C(_1225__bF_buf5), .Y(_1218__22_) );
	OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag1_23_), .Y(_1271_) );
	NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_21_), .B(_1249__bF_buf0), .Y(_1272_) );
	AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1271_), .C(_1225__bF_buf4), .Y(_1218__23_) );
	OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag1_24_), .Y(_1273_) );
	NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_22_), .B(_1249__bF_buf3), .Y(_1274_) );
	AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1273_), .C(_1225__bF_buf3), .Y(_1218__24_) );
	OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag1_25_), .Y(_1275_) );
	NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_23_), .B(_1249__bF_buf2), .Y(_1276_) );
	AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1275_), .C(_1225__bF_buf2), .Y(_1218__25_) );
	OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag1_26_), .Y(_1277_) );
	NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_24_), .B(_1249__bF_buf1), .Y(_1278_) );
	AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1277_), .C(_1225__bF_buf1), .Y(_1218__26_) );
	OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag1_27_), .Y(_1279_) );
	NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_25_), .B(_1249__bF_buf0), .Y(_1280_) );
	AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1279_), .C(_1225__bF_buf0), .Y(_1218__27_) );
	OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag1_28_), .Y(_1281_) );
	NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_26_), .B(_1249__bF_buf3), .Y(_1282_) );
	AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1281_), .C(_1225__bF_buf5), .Y(_1218__28_) );
	OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag1_29_), .Y(_1283_) );
	NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_27_), .B(_1249__bF_buf2), .Y(_1284_) );
	AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1283_), .C(_1225__bF_buf4), .Y(_1218__29_) );
	OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag1_30_), .Y(_1285_) );
	NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_28_), .B(_1249__bF_buf1), .Y(_1286_) );
	AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1285_), .C(_1225__bF_buf3), .Y(_1218__30_) );
	OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag1_31_), .Y(_1287_) );
	NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_29_), .B(_1249__bF_buf0), .Y(_1288_) );
	AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1288_), .B(_1287_), .C(_1225__bF_buf2), .Y(_1218__31_) );
	OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag1_32_), .Y(_1289_) );
	NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_30_), .B(_1249__bF_buf3), .Y(_1290_) );
	AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1289_), .C(_1225__bF_buf1), .Y(_1218__32_) );
	OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag1_33_), .Y(_1291_) );
	NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_31_), .B(_1249__bF_buf2), .Y(_1292_) );
	AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1291_), .C(_1225__bF_buf0), .Y(_1218__33_) );
	INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_0_), .Y(_1293_) );
	OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_0_), .B(_1228__bF_buf2), .C(_1224__bF_buf0), .Y(_1294_) );
	AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1228__bF_buf1), .C(_1294_), .Y(_1219__0_) );
	INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_1_), .Y(_1295_) );
	OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_1_), .B(_1228__bF_buf0), .C(_1224__bF_buf3), .Y(_1296_) );
	AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1228__bF_buf5), .C(_1296_), .Y(_1219__1_) );
	INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_2_), .Y(_1297_) );
	OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_2_), .B(_1228__bF_buf4), .C(_1224__bF_buf2), .Y(_1298_) );
	AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .B(_1228__bF_buf3), .C(_1298_), .Y(_1219__2_) );
	INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_3_), .Y(_1299_) );
	OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_3_), .B(_1228__bF_buf2), .C(_1224__bF_buf1), .Y(_1300_) );
	AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1228__bF_buf1), .C(_1300_), .Y(_1219__3_) );
	INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_4_), .Y(_1301_) );
	OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_4_), .B(_1228__bF_buf0), .C(_1224__bF_buf0), .Y(_1302_) );
	AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1301_), .B(_1228__bF_buf5), .C(_1302_), .Y(_1219__4_) );
	INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_5_), .Y(_1303_) );
	OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_5_), .B(_1228__bF_buf4), .C(_1224__bF_buf3), .Y(_1304_) );
	AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1228__bF_buf3), .C(_1304_), .Y(_1219__5_) );
	INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_6_), .Y(_1305_) );
	OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_6_), .B(_1228__bF_buf2), .C(_1224__bF_buf2), .Y(_1306_) );
	AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_1228__bF_buf1), .C(_1306_), .Y(_1219__6_) );
	INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_7_), .Y(_1307_) );
	OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_7_), .B(_1228__bF_buf0), .C(_1224__bF_buf1), .Y(_1308_) );
	AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1228__bF_buf5), .C(_1308_), .Y(_1219__7_) );
	INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_8_), .Y(_1309_) );
	OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_8_), .B(_1228__bF_buf4), .C(_1224__bF_buf0), .Y(_1310_) );
	AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1228__bF_buf3), .C(_1310_), .Y(_1219__8_) );
	INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_9_), .Y(_1311_) );
	OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_9_), .B(_1228__bF_buf2), .C(_1224__bF_buf3), .Y(_1312_) );
	AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1228__bF_buf1), .C(_1312_), .Y(_1219__9_) );
	INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_10_), .Y(_1313_) );
	OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_10_), .B(_1228__bF_buf0), .C(_1224__bF_buf2), .Y(_1314_) );
	AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1228__bF_buf5), .C(_1314_), .Y(_1219__10_) );
	INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_11_), .Y(_1315_) );
	OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_11_), .B(_1228__bF_buf4), .C(_1224__bF_buf1), .Y(_1316_) );
	AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .B(_1228__bF_buf3), .C(_1316_), .Y(_1219__11_) );
	OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag2_12_), .Y(_1317_) );
	AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1317_), .C(_1225__bF_buf5), .Y(_1219__12_) );
	OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag2_13_), .Y(_1318_) );
	AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1318_), .C(_1225__bF_buf4), .Y(_1219__13_) );
	OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag2_14_), .Y(_1319_) );
	AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1319_), .C(_1225__bF_buf3), .Y(_1219__14_) );
	OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag2_15_), .Y(_1320_) );
	AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1320_), .C(_1225__bF_buf2), .Y(_1219__15_) );
	OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag2_16_), .Y(_1321_) );
	AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_1321_), .C(_1225__bF_buf1), .Y(_1219__16_) );
	OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag2_17_), .Y(_1322_) );
	AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1322_), .C(_1225__bF_buf0), .Y(_1219__17_) );
	OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag2_18_), .Y(_1323_) );
	AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1323_), .C(_1225__bF_buf5), .Y(_1219__18_) );
	OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag2_19_), .Y(_1324_) );
	AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1324_), .C(_1225__bF_buf4), .Y(_1219__19_) );
	OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag2_20_), .Y(_1325_) );
	AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1325_), .C(_1225__bF_buf3), .Y(_1219__20_) );
	OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag2_21_), .Y(_1326_) );
	AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1326_), .C(_1225__bF_buf2), .Y(_1219__21_) );
	OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag2_22_), .Y(_1327_) );
	AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1327_), .C(_1225__bF_buf1), .Y(_1219__22_) );
	OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag2_23_), .Y(_1328_) );
	AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1328_), .C(_1225__bF_buf0), .Y(_1219__23_) );
	OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag2_24_), .Y(_1329_) );
	AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1329_), .C(_1225__bF_buf5), .Y(_1219__24_) );
	OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag2_25_), .Y(_1330_) );
	AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1330_), .C(_1225__bF_buf4), .Y(_1219__25_) );
	OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag2_26_), .Y(_1331_) );
	AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1331_), .C(_1225__bF_buf3), .Y(_1219__26_) );
	OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag2_27_), .Y(_1332_) );
	AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1332_), .C(_1225__bF_buf2), .Y(_1219__27_) );
	OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1222__bF_buf1), .C(biu_mmu_reg_ag2_28_), .Y(_1333_) );
	AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1333_), .C(_1225__bF_buf1), .Y(_1219__28_) );
	OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf5), .B(_1222__bF_buf0), .C(biu_mmu_reg_ag2_29_), .Y(_1334_) );
	AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1334_), .C(_1225__bF_buf0), .Y(_1219__29_) );
	OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf4), .B(_1222__bF_buf5), .C(biu_mmu_reg_ag2_30_), .Y(_1335_) );
	AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1335_), .C(_1225__bF_buf5), .Y(_1219__30_) );
	OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf3), .B(_1222__bF_buf4), .C(biu_mmu_reg_ag2_31_), .Y(_1336_) );
	AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1288_), .B(_1336_), .C(_1225__bF_buf4), .Y(_1219__31_) );
	OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf2), .B(_1222__bF_buf3), .C(biu_mmu_reg_ag2_32_), .Y(_1337_) );
	AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1337_), .C(_1225__bF_buf3), .Y(_1219__32_) );
	OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf1), .B(_1222__bF_buf2), .C(biu_mmu_reg_ag2_33_), .Y(_1338_) );
	AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1338_), .C(_1225__bF_buf2), .Y(_1219__33_) );
	INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_3_), .Y(_1339_) );
	INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf2), .Y(_1340_) );
	NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_exce_chk_statu_biu_6_bF_buf1), .Y(_1341_) );
	AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1340_), .C(_1339_), .Y(_1342_) );
	NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1340_), .C(_1341_), .Y(_1343_) );
	INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .Y(_1344_) );
	NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1344_), .Y(biu_mmu_pte_new_7_) );
	AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_0_), .Y(biu_mmu_pte_new_0_) );
	AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_1_), .Y(biu_mmu_pte_new_1_) );
	AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_2_), .Y(biu_mmu_pte_new_2_) );
	AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_3_), .Y(biu_mmu_pte_new_3_) );
	AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_4_), .Y(biu_mmu_pte_new_4_) );
	AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_5_), .Y(biu_mmu_pte_new_5_) );
	AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_8_), .Y(biu_mmu_pte_new_8_) );
	AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_9_), .Y(biu_mmu_pte_new_9_) );
	AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_10_), .Y(biu_mmu_pte_new_10_) );
	AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_11_), .Y(biu_mmu_pte_new_11_) );
	AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_12_), .Y(biu_mmu_pte_new_12_) );
	AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_13_), .Y(biu_mmu_pte_new_13_) );
	AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_14_), .Y(biu_mmu_pte_new_14_) );
	AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_15_), .Y(biu_mmu_pte_new_15_) );
	AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_16_), .Y(biu_mmu_pte_new_16_) );
	AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_17_), .Y(biu_mmu_pte_new_17_) );
	AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_18_), .Y(biu_mmu_pte_new_18_) );
	AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_19_), .Y(biu_mmu_pte_new_19_) );
	AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_20_), .Y(biu_mmu_pte_new_20_) );
	AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_21_), .Y(biu_mmu_pte_new_21_) );
	AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_22_), .Y(biu_mmu_pte_new_22_) );
	AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_23_), .Y(biu_mmu_pte_new_23_) );
	AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_24_), .Y(biu_mmu_pte_new_24_) );
	AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_25_), .Y(biu_mmu_pte_new_25_) );
	AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_26_), .Y(biu_mmu_pte_new_26_) );
	AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf2), .B(biu_ahb_data_out_27_), .Y(biu_mmu_pte_new_27_) );
	AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf1), .B(biu_ahb_data_out_28_), .Y(biu_mmu_pte_new_28_) );
	AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf0), .B(biu_ahb_data_out_29_), .Y(biu_mmu_pte_new_29_) );
	AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf4), .B(biu_ahb_data_out_30_), .Y(biu_mmu_pte_new_30_) );
	AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_pte_new_7_bF_buf3), .B(biu_ahb_data_out_31_), .Y(biu_mmu_pte_new_31_) );
	NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1341_), .Y(_1345_) );
	OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf1), .B(biu_exce_chk_statu_biu_5_), .C(biu_exce_chk_statu_biu_6_bF_buf0), .Y(_1346_) );
	NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_0_), .B(_1339_), .Y(_1347_) );
	NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .B(_1347_), .Y(_1348_) );
	NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1346_), .C(_1348_), .Y(_1349_) );
	INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_sum), .Y(_1350_) );
	INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .Y(_1351_) );
	NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf4), .B(_1351_), .Y(_1352_) );
	OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1352_), .C(biu_ahb_data_out_4_), .Y(_1353_) );
	INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_1_), .Y(_1354_) );
	NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_mxr), .B(_1354_), .Y(_1355_) );
	NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_3_), .B(_1341_), .Y(_1356_) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .B(biu_exce_chk_statu_biu_6_bF_buf3), .Y(_1357_) );
	INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_3_), .Y(_1358_) );
	NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf0), .B(_1358_), .Y(_1359_) );
	OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_7_), .B(biu_ahb_data_out_6_), .C(biu_ahb_data_out_0_), .Y(_1360_) );
	INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .Y(_1361_) );
	OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1359_), .C(_1361_), .Y(_1362_) );
	AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1356_), .C(_1362_), .Y(_1363_) );
	AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1353_), .C(_1349_), .Y(biu_exce_chk_mmu_ld_page_fault) );
	INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_0_), .Y(_1364_) );
	INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_2_), .Y(_1365_) );
	NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(_1365_), .Y(_1366_) );
	NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1220__bF_buf0), .B(_1366_), .Y(_1367_) );
	NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_0_), .B(_1228__bF_buf2), .Y(_1368_) );
	AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1367_), .C(_1343_), .D(_1368_), .Y(_1369_) );
	INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_5_), .Y(_1370_) );
	OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1370_), .C(_1346_), .Y(_1371_) );
	NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_2_), .B(_1347_), .C(_1366_), .Y(_1372_) );
	NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_7_), .B(biu_ahb_data_out_6_), .Y(_1373_) );
	AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(biu_ahb_data_out_4_), .Y(_1374_) );
	AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1374_), .C(_1371_), .D(_1372_), .Y(_1375_) );
	NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1375_), .Y(biu_exce_chk_mmu_st_page_fault) );
	OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_4_bF_buf3), .B(_1357_), .C(_1348_), .Y(_1376_) );
	NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(biu_ahb_data_out_0_), .B(_1376_), .Y(biu_exce_chk_page_not_value) );
	INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .Y(_1377_) );
	NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_0_), .B(_1377__bF_buf3), .Y(_1378_) );
	NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_biu_1_), .B(_1365_), .Y(_1379_) );
	INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(_1379__bF_buf4), .Y(_1380_) );
	OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1380_), .C(_1378_), .Y(biu_addr_mmu_0_) );
	NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_1_), .B(_1377__bF_buf2), .Y(_1381_) );
	OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1380_), .C(_1381_), .Y(biu_addr_mmu_1_) );
	AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_22_), .B(_1221__bF_buf1), .C(biu_mmu_reg_ag2_2_), .D(_1379__bF_buf3), .Y(_1382_) );
	OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .B(_1366_), .C(_1382_), .Y(biu_addr_mmu_2_) );
	AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_23_), .B(_1221__bF_buf0), .C(biu_mmu_reg_ag2_3_), .D(_1379__bF_buf2), .Y(_1383_) );
	OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1366_), .C(_1383_), .Y(biu_addr_mmu_3_) );
	AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_24_), .B(_1221__bF_buf4), .C(biu_mmu_reg_ag2_4_), .D(_1379__bF_buf1), .Y(_1384_) );
	OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1366_), .C(_1384_), .Y(biu_addr_mmu_4_) );
	AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_25_), .B(_1221__bF_buf3), .C(biu_mmu_reg_ag2_5_), .D(_1379__bF_buf0), .Y(_1385_) );
	OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1366_), .C(_1385_), .Y(biu_addr_mmu_5_) );
	AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_26_), .B(_1221__bF_buf2), .C(biu_mmu_reg_ag2_6_), .D(_1379__bF_buf4), .Y(_1386_) );
	OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1366_), .C(_1386_), .Y(biu_addr_mmu_6_) );
	AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_27_), .B(_1221__bF_buf1), .C(biu_mmu_reg_ag2_7_), .D(_1379__bF_buf3), .Y(_1387_) );
	OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1366_), .C(_1387_), .Y(biu_addr_mmu_7_) );
	AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_28_), .B(_1221__bF_buf0), .C(biu_mmu_reg_ag2_8_), .D(_1379__bF_buf2), .Y(_1388_) );
	OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_1366_), .C(_1388_), .Y(biu_addr_mmu_8_) );
	AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_29_), .B(_1221__bF_buf4), .C(biu_mmu_reg_ag2_9_), .D(_1379__bF_buf1), .Y(_1389_) );
	OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_1366_), .C(_1389_), .Y(biu_addr_mmu_9_) );
	AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_30_), .B(_1221__bF_buf3), .C(biu_mmu_reg_ag2_10_), .D(_1379__bF_buf0), .Y(_1390_) );
	OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1366_), .C(_1390_), .Y(biu_addr_mmu_10_) );
	AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(biu_addr_mmu_in_31_), .B(_1221__bF_buf2), .C(biu_mmu_reg_ag2_11_), .D(_1379__bF_buf4), .Y(_1391_) );
	OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1366_), .C(_1391_), .Y(biu_addr_mmu_11_) );
	NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_12_), .B(_1377__bF_buf1), .Y(_1392_) );
	NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_12_), .B(_1379__bF_buf3), .Y(_1393_) );
	NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_12_), .B(_1221__bF_buf1), .Y(_1394_) );
	NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1394_), .C(_1392_), .Y(biu_addr_mmu_12_) );
	NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_13_), .B(_1377__bF_buf0), .Y(_1395_) );
	NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_13_), .B(_1379__bF_buf2), .Y(_1396_) );
	NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_13_), .B(_1221__bF_buf0), .Y(_1397_) );
	NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1396_), .B(_1397_), .C(_1395_), .Y(biu_addr_mmu_13_) );
	NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_14_), .B(_1377__bF_buf3), .Y(_1398_) );
	NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_14_), .B(_1379__bF_buf1), .Y(_1399_) );
	NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_14_), .B(_1221__bF_buf4), .Y(_1400_) );
	NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1400_), .C(_1398_), .Y(biu_addr_mmu_14_) );
	NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_15_), .B(_1377__bF_buf2), .Y(_1401_) );
	NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_15_), .B(_1379__bF_buf0), .Y(_1402_) );
	NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_15_), .B(_1221__bF_buf3), .Y(_1403_) );
	NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1403_), .C(_1401_), .Y(biu_addr_mmu_15_) );
	NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_16_), .B(_1377__bF_buf1), .Y(_1404_) );
	NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_16_), .B(_1379__bF_buf4), .Y(_1405_) );
	NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_16_), .B(_1221__bF_buf2), .Y(_1406_) );
	NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1406_), .C(_1404_), .Y(biu_addr_mmu_16_) );
	NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_17_), .B(_1377__bF_buf0), .Y(_1407_) );
	NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_17_), .B(_1379__bF_buf3), .Y(_1408_) );
	NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_17_), .B(_1221__bF_buf1), .Y(_1409_) );
	NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1409_), .C(_1407_), .Y(biu_addr_mmu_17_) );
	NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_18_), .B(_1377__bF_buf3), .Y(_1410_) );
	NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_18_), .B(_1379__bF_buf2), .Y(_1411_) );
	NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_18_), .B(_1221__bF_buf0), .Y(_1412_) );
	NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1412_), .C(_1410_), .Y(biu_addr_mmu_18_) );
	NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_19_), .B(_1377__bF_buf2), .Y(_1413_) );
	NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_19_), .B(_1379__bF_buf1), .Y(_1414_) );
	NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_19_), .B(_1221__bF_buf4), .Y(_1415_) );
	NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1415_), .C(_1413_), .Y(biu_addr_mmu_19_) );
	NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_20_), .B(_1377__bF_buf1), .Y(_1416_) );
	NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_20_), .B(_1379__bF_buf0), .Y(_1417_) );
	NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_20_), .B(_1221__bF_buf3), .Y(_1418_) );
	NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1418_), .C(_1416_), .Y(biu_addr_mmu_20_) );
	NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_21_), .B(_1377__bF_buf0), .Y(_1419_) );
	NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_21_), .B(_1379__bF_buf4), .Y(_1420_) );
	NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_21_), .B(_1221__bF_buf2), .Y(_1421_) );
	NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1421_), .C(_1419_), .Y(biu_addr_mmu_21_) );
	NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_22_), .B(_1377__bF_buf3), .Y(_1422_) );
	NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_22_), .B(_1379__bF_buf3), .Y(_1423_) );
	NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_22_), .B(_1221__bF_buf1), .Y(_1424_) );
	NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1423_), .B(_1424_), .C(_1422_), .Y(biu_addr_mmu_22_) );
	NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_23_), .B(_1377__bF_buf2), .Y(_1425_) );
	NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_23_), .B(_1379__bF_buf2), .Y(_1426_) );
	NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_23_), .B(_1221__bF_buf0), .Y(_1427_) );
	NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1427_), .C(_1425_), .Y(biu_addr_mmu_23_) );
	NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_24_), .B(_1377__bF_buf1), .Y(_1428_) );
	NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_24_), .B(_1379__bF_buf1), .Y(_1429_) );
	NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_24_), .B(_1221__bF_buf4), .Y(_1430_) );
	NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1429_), .B(_1430_), .C(_1428_), .Y(biu_addr_mmu_24_) );
	NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_25_), .B(_1377__bF_buf0), .Y(_1431_) );
	NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_25_), .B(_1379__bF_buf0), .Y(_1432_) );
	NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_25_), .B(_1221__bF_buf3), .Y(_1433_) );
	NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1433_), .C(_1431_), .Y(biu_addr_mmu_25_) );
	NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_26_), .B(_1377__bF_buf3), .Y(_1434_) );
	NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_26_), .B(_1379__bF_buf4), .Y(_1435_) );
	NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_26_), .B(_1221__bF_buf2), .Y(_1436_) );
	NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_1436_), .C(_1434_), .Y(biu_addr_mmu_26_) );
	NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_27_), .B(_1377__bF_buf2), .Y(_1437_) );
	NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_27_), .B(_1379__bF_buf3), .Y(_1438_) );
	NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_27_), .B(_1221__bF_buf1), .Y(_1439_) );
	NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1439_), .C(_1437_), .Y(biu_addr_mmu_27_) );
	NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_28_), .B(_1377__bF_buf1), .Y(_1440_) );
	NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_28_), .B(_1379__bF_buf2), .Y(_1441_) );
	NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_28_), .B(_1221__bF_buf0), .Y(_1442_) );
	NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1442_), .C(_1440_), .Y(biu_addr_mmu_28_) );
	NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_29_), .B(_1377__bF_buf0), .Y(_1443_) );
	NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_29_), .B(_1379__bF_buf1), .Y(_1444_) );
	NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_29_), .B(_1221__bF_buf4), .Y(_1445_) );
	NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .B(_1445_), .C(_1443_), .Y(biu_addr_mmu_29_) );
	NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_30_), .B(_1377__bF_buf3), .Y(_1446_) );
	NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_30_), .B(_1379__bF_buf0), .Y(_1447_) );
	NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_30_), .B(_1221__bF_buf3), .Y(_1448_) );
	NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1448_), .C(_1446_), .Y(biu_addr_mmu_30_) );
	NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_31_), .B(_1377__bF_buf2), .Y(_1449_) );
	NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_31_), .B(_1379__bF_buf4), .Y(_1450_) );
	NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_31_), .B(_1221__bF_buf2), .Y(_1451_) );
	NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1451_), .C(_1449_), .Y(biu_addr_mmu_31_) );
	NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_32_), .B(_1377__bF_buf1), .Y(_1452_) );
	NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_32_), .B(_1379__bF_buf3), .Y(_1453_) );
	NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_32_), .B(_1221__bF_buf1), .Y(_1454_) );
	NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1454_), .C(_1452_), .Y(biu_addr_mmu_32_) );
	NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag1_33_), .B(_1377__bF_buf0), .Y(_1455_) );
	NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_reg_ag2_33_), .B(_1379__bF_buf2), .Y(_1456_) );
	NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_33_), .B(_1221__bF_buf0), .Y(_1457_) );
	NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(_1457_), .C(_1455_), .Y(biu_addr_mmu_33_) );
	DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1218__0_), .Q(biu_mmu_reg_ag1_0_) );
	DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_1218__1_), .Q(biu_mmu_reg_ag1_1_) );
	DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_1218__2_), .Q(biu_mmu_reg_ag1_2_) );
	DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_1218__3_), .Q(biu_mmu_reg_ag1_3_) );
	DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1218__4_), .Q(biu_mmu_reg_ag1_4_) );
	DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_1218__5_), .Q(biu_mmu_reg_ag1_5_) );
	DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_1218__6_), .Q(biu_mmu_reg_ag1_6_) );
	DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_1218__7_), .Q(biu_mmu_reg_ag1_7_) );
	DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_1218__8_), .Q(biu_mmu_reg_ag1_8_) );
	DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_1218__9_), .Q(biu_mmu_reg_ag1_9_) );
	DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_1218__10_), .Q(biu_mmu_reg_ag1_10_) );
	DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_1218__11_), .Q(biu_mmu_reg_ag1_11_) );
	DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_1218__12_), .Q(biu_mmu_reg_ag1_12_) );
	DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_1218__13_), .Q(biu_mmu_reg_ag1_13_) );
	DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_1218__14_), .Q(biu_mmu_reg_ag1_14_) );
	DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_1218__15_), .Q(biu_mmu_reg_ag1_15_) );
	DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_1218__16_), .Q(biu_mmu_reg_ag1_16_) );
	DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_1218__17_), .Q(biu_mmu_reg_ag1_17_) );
	DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_1218__18_), .Q(biu_mmu_reg_ag1_18_) );
	DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_1218__19_), .Q(biu_mmu_reg_ag1_19_) );
	DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_1218__20_), .Q(biu_mmu_reg_ag1_20_) );
	DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_1218__21_), .Q(biu_mmu_reg_ag1_21_) );
	DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_1218__22_), .Q(biu_mmu_reg_ag1_22_) );
	DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_1218__23_), .Q(biu_mmu_reg_ag1_23_) );
	DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_1218__24_), .Q(biu_mmu_reg_ag1_24_) );
	DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_1218__25_), .Q(biu_mmu_reg_ag1_25_) );
	DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_1218__26_), .Q(biu_mmu_reg_ag1_26_) );
	DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_1218__27_), .Q(biu_mmu_reg_ag1_27_) );
	DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_1218__28_), .Q(biu_mmu_reg_ag1_28_) );
	DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1218__29_), .Q(biu_mmu_reg_ag1_29_) );
	DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_1218__30_), .Q(biu_mmu_reg_ag1_30_) );
	DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_1218__31_), .Q(biu_mmu_reg_ag1_31_) );
	DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_1218__32_), .Q(biu_mmu_reg_ag1_32_) );
	DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_1218__33_), .Q(biu_mmu_reg_ag1_33_) );
	DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_1219__0_), .Q(biu_mmu_reg_ag2_0_) );
	DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_1219__1_), .Q(biu_mmu_reg_ag2_1_) );
	DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1219__2_), .Q(biu_mmu_reg_ag2_2_) );
	DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_1219__3_), .Q(biu_mmu_reg_ag2_3_) );
	DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_1219__4_), .Q(biu_mmu_reg_ag2_4_) );
	DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_1219__5_), .Q(biu_mmu_reg_ag2_5_) );
	DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_1219__6_), .Q(biu_mmu_reg_ag2_6_) );
	DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_1219__7_), .Q(biu_mmu_reg_ag2_7_) );
	DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_1219__8_), .Q(biu_mmu_reg_ag2_8_) );
	DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_1219__9_), .Q(biu_mmu_reg_ag2_9_) );
	DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_1219__10_), .Q(biu_mmu_reg_ag2_10_) );
	DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1219__11_), .Q(biu_mmu_reg_ag2_11_) );
	DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1219__12_), .Q(biu_mmu_reg_ag2_12_) );
	DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1219__13_), .Q(biu_mmu_reg_ag2_13_) );
	DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1219__14_), .Q(biu_mmu_reg_ag2_14_) );
	DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1219__15_), .Q(biu_mmu_reg_ag2_15_) );
	DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1219__16_), .Q(biu_mmu_reg_ag2_16_) );
	DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1219__17_), .Q(biu_mmu_reg_ag2_17_) );
	DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1219__18_), .Q(biu_mmu_reg_ag2_18_) );
	DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1219__19_), .Q(biu_mmu_reg_ag2_19_) );
	DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1219__20_), .Q(biu_mmu_reg_ag2_20_) );
	DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1219__21_), .Q(biu_mmu_reg_ag2_21_) );
	DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1219__22_), .Q(biu_mmu_reg_ag2_22_) );
	DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_1219__23_), .Q(biu_mmu_reg_ag2_23_) );
	DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_1219__24_), .Q(biu_mmu_reg_ag2_24_) );
	DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_1219__25_), .Q(biu_mmu_reg_ag2_25_) );
	DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_1219__26_), .Q(biu_mmu_reg_ag2_26_) );
	DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_1219__27_), .Q(biu_mmu_reg_ag2_27_) );
	DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_1219__28_), .Q(biu_mmu_reg_ag2_28_) );
	DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_1219__29_), .Q(biu_mmu_reg_ag2_29_) );
	DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_1219__30_), .Q(biu_mmu_reg_ag2_30_) );
	DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_1219__31_), .Q(biu_mmu_reg_ag2_31_) );
	DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_1219__32_), .Q(biu_mmu_reg_ag2_32_) );
	DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_1219__33_), .Q(biu_mmu_reg_ag2_33_) );
	INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .Y(_2460_) );
	NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(biu_ins_7_), .Y(_2461_) );
	NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_9_), .B(biu_ins_10_), .Y(_2462_) );
	NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2462_), .Y(_2463_) );
	NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .B(_2463_), .Y(_2464_) );
	NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_2_), .Y(_2465_) );
	NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(biu_exce_chk_statu_cpu_0_), .Y(_2466_) );
	INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .Y(_2467_) );
	NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_wr), .B(_2465_), .C(_2467_), .Y(_2468_) );
	NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_2468_), .B(_2464_), .Y(_2469_) );
	INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_7_), .Y(_2470_) );
	NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(_2470_), .Y(_2471_) );
	INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .Y(_2472_) );
	AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2472_), .Y(_2473_) );
	INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .Y(_2474_) );
	AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2462_), .C(_2474_), .Y(_2475_) );
	NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2464_), .Y(_2476_) );
	INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_9_), .Y(_2477_) );
	NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2461_), .Y(_2478_) );
	NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_10_), .B(_2478_), .Y(_2479_) );
	AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2479_), .C(_2476_), .Y(_2480_) );
	OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(biu_ins_7_), .C(biu_ins_9_), .Y(_2481_) );
	NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2481_), .B(_2478_), .Y(_2482_) );
	NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2480_), .C(_2473__bF_buf7), .Y(_2483_) );
	NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(_2470_), .C(_2469_), .Y(_2484_) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2475_), .Y(_2485_) );
	NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2479_), .Y(_2486_) );
	NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2486_), .C(_2485_), .Y(_2487_) );
	OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_29__0_), .Y(_2488_) );
	OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf4), .B(_2483__bF_buf4), .C(_2488_), .Y(_2332_) );
	INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .Y(_2489_) );
	OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_29__1_), .Y(_2490_) );
	OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf4), .B(_2483__bF_buf3), .C(_2490_), .Y(_2333_) );
	INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .Y(_2491_) );
	OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_29__2_), .Y(_2492_) );
	OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf4), .B(_2483__bF_buf2), .C(_2492_), .Y(_2334_) );
	INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .Y(_2493_) );
	OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_29__3_), .Y(_2494_) );
	OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf4), .B(_2483__bF_buf1), .C(_2494_), .Y(_2335_) );
	INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .Y(_2495_) );
	OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_29__4_), .Y(_2496_) );
	OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf4), .B(_2483__bF_buf0), .C(_2496_), .Y(_2336_) );
	INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .Y(_2497_) );
	OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_29__5_), .Y(_2498_) );
	OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf4), .B(_2483__bF_buf4), .C(_2498_), .Y(_2337_) );
	INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .Y(_2499_) );
	OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_29__6_), .Y(_2500_) );
	OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf4), .B(_2483__bF_buf3), .C(_2500_), .Y(_2338_) );
	INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .Y(_2501_) );
	OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_29__7_), .Y(_2502_) );
	OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf4), .B(_2483__bF_buf2), .C(_2502_), .Y(_2339_) );
	INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .Y(_2503_) );
	OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_29__8_), .Y(_2504_) );
	OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf4), .B(_2483__bF_buf1), .C(_2504_), .Y(_2340_) );
	INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .Y(_2505_) );
	OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_29__9_), .Y(_2506_) );
	OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf4), .B(_2483__bF_buf0), .C(_2506_), .Y(_2341_) );
	INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .Y(_2507_) );
	OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_29__10_), .Y(_2508_) );
	OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf4), .B(_2483__bF_buf4), .C(_2508_), .Y(_2342_) );
	INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .Y(_2509_) );
	OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_29__11_), .Y(_2510_) );
	OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf4), .B(_2483__bF_buf3), .C(_2510_), .Y(_2343_) );
	INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .Y(_2511_) );
	OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_29__12_), .Y(_2512_) );
	OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf4), .B(_2483__bF_buf2), .C(_2512_), .Y(_2344_) );
	INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .Y(_2513_) );
	OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_29__13_), .Y(_2514_) );
	OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf4), .B(_2483__bF_buf1), .C(_2514_), .Y(_2345_) );
	INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .Y(_2515_) );
	OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_29__14_), .Y(_2516_) );
	OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf4), .B(_2483__bF_buf0), .C(_2516_), .Y(_2346_) );
	INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .Y(_2517_) );
	OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_29__15_), .Y(_2518_) );
	OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf4), .B(_2483__bF_buf4), .C(_2518_), .Y(_2347_) );
	INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .Y(_2519_) );
	OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_29__16_), .Y(_2520_) );
	OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf4), .B(_2483__bF_buf3), .C(_2520_), .Y(_2348_) );
	INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .Y(_2521_) );
	OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_29__17_), .Y(_2522_) );
	OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf4), .B(_2483__bF_buf2), .C(_2522_), .Y(_2349_) );
	INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .Y(_2523_) );
	OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_29__18_), .Y(_2524_) );
	OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf4), .B(_2483__bF_buf1), .C(_2524_), .Y(_2350_) );
	INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .Y(_2525_) );
	OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_29__19_), .Y(_2526_) );
	OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf4), .B(_2483__bF_buf0), .C(_2526_), .Y(_2351_) );
	INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .Y(_2527_) );
	OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_29__20_), .Y(_2528_) );
	OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf4), .B(_2483__bF_buf4), .C(_2528_), .Y(_2352_) );
	INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .Y(_2529_) );
	OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_29__21_), .Y(_2530_) );
	OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf4), .B(_2483__bF_buf3), .C(_2530_), .Y(_2353_) );
	INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .Y(_2531_) );
	OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_29__22_), .Y(_2532_) );
	OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf4), .B(_2483__bF_buf2), .C(_2532_), .Y(_2354_) );
	INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .Y(_2533_) );
	OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_29__23_), .Y(_2534_) );
	OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf4), .B(_2483__bF_buf1), .C(_2534_), .Y(_2355_) );
	INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .Y(_2535_) );
	OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_29__24_), .Y(_2536_) );
	OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf4), .B(_2483__bF_buf0), .C(_2536_), .Y(_2356_) );
	INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .Y(_2537_) );
	OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_29__25_), .Y(_2538_) );
	OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf4), .B(_2483__bF_buf4), .C(_2538_), .Y(_2357_) );
	INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .Y(_2539_) );
	OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_29__26_), .Y(_2540_) );
	OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf4), .B(_2483__bF_buf3), .C(_2540_), .Y(_2358_) );
	INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .Y(_2541_) );
	OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_29__27_), .Y(_2542_) );
	OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf4), .B(_2483__bF_buf2), .C(_2542_), .Y(_2359_) );
	INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .Y(_2543_) );
	OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_29__28_), .Y(_2544_) );
	OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf4), .B(_2483__bF_buf1), .C(_2544_), .Y(_2360_) );
	INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .Y(_2545_) );
	OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_29__29_), .Y(_2546_) );
	OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf4), .B(_2483__bF_buf0), .C(_2546_), .Y(_2361_) );
	INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .Y(_2547_) );
	OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_29__30_), .Y(_2548_) );
	OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_2483__bF_buf4), .C(_2548_), .Y(_2362_) );
	INVX8 INVX8_44 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .Y(_2549_) );
	OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_29__31_), .Y(_2550_) );
	OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf4), .B(_2483__bF_buf3), .C(_2550_), .Y(_2363_) );
	INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .Y(_2551_) );
	NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2480_), .C(_2473__bF_buf6), .Y(_2552_) );
	NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2486_), .C(_2485_), .Y(_2553_) );
	OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_25__0_), .Y(_2554_) );
	OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf3), .B(_2552__bF_buf4), .C(_2554_), .Y(_2364_) );
	OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_25__1_), .Y(_2555_) );
	OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf3), .B(_2552__bF_buf3), .C(_2555_), .Y(_2365_) );
	OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_25__2_), .Y(_2556_) );
	OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf3), .B(_2552__bF_buf2), .C(_2556_), .Y(_2366_) );
	OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_25__3_), .Y(_2557_) );
	OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf3), .B(_2552__bF_buf1), .C(_2557_), .Y(_2367_) );
	OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_25__4_), .Y(_2558_) );
	OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf3), .B(_2552__bF_buf0), .C(_2558_), .Y(_2368_) );
	OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_25__5_), .Y(_2559_) );
	OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf3), .B(_2552__bF_buf4), .C(_2559_), .Y(_2369_) );
	OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_25__6_), .Y(_2560_) );
	OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf3), .B(_2552__bF_buf3), .C(_2560_), .Y(_2370_) );
	OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_25__7_), .Y(_2561_) );
	OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf3), .B(_2552__bF_buf2), .C(_2561_), .Y(_2371_) );
	OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_25__8_), .Y(_2562_) );
	OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf3), .B(_2552__bF_buf1), .C(_2562_), .Y(_2372_) );
	OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_25__9_), .Y(_2563_) );
	OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf3), .B(_2552__bF_buf0), .C(_2563_), .Y(_2373_) );
	OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_25__10_), .Y(_2564_) );
	OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf3), .B(_2552__bF_buf4), .C(_2564_), .Y(_2374_) );
	OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_25__11_), .Y(_2565_) );
	OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf3), .B(_2552__bF_buf3), .C(_2565_), .Y(_2375_) );
	OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_25__12_), .Y(_2566_) );
	OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf3), .B(_2552__bF_buf2), .C(_2566_), .Y(_2376_) );
	OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_25__13_), .Y(_2567_) );
	OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf3), .B(_2552__bF_buf1), .C(_2567_), .Y(_2377_) );
	OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_25__14_), .Y(_2568_) );
	OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf3), .B(_2552__bF_buf0), .C(_2568_), .Y(_2378_) );
	OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_25__15_), .Y(_2569_) );
	OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf3), .B(_2552__bF_buf4), .C(_2569_), .Y(_2379_) );
	OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_25__16_), .Y(_2570_) );
	OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf3), .B(_2552__bF_buf3), .C(_2570_), .Y(_2380_) );
	OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_25__17_), .Y(_2571_) );
	OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf3), .B(_2552__bF_buf2), .C(_2571_), .Y(_2381_) );
	OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_25__18_), .Y(_2572_) );
	OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf3), .B(_2552__bF_buf1), .C(_2572_), .Y(_2382_) );
	OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_25__19_), .Y(_2573_) );
	OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf3), .B(_2552__bF_buf0), .C(_2573_), .Y(_2383_) );
	OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_25__20_), .Y(_2574_) );
	OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf3), .B(_2552__bF_buf4), .C(_2574_), .Y(_2384_) );
	OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_25__21_), .Y(_2575_) );
	OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf3), .B(_2552__bF_buf3), .C(_2575_), .Y(_2385_) );
	OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_25__22_), .Y(_2576_) );
	OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf3), .B(_2552__bF_buf2), .C(_2576_), .Y(_2386_) );
	OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_25__23_), .Y(_2577_) );
	OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf3), .B(_2552__bF_buf1), .C(_2577_), .Y(_2387_) );
	OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_25__24_), .Y(_2578_) );
	OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf3), .B(_2552__bF_buf0), .C(_2578_), .Y(_2388_) );
	OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_25__25_), .Y(_2579_) );
	OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf3), .B(_2552__bF_buf4), .C(_2579_), .Y(_2389_) );
	OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_25__26_), .Y(_2580_) );
	OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf3), .B(_2552__bF_buf3), .C(_2580_), .Y(_2390_) );
	OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_25__27_), .Y(_2581_) );
	OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf3), .B(_2552__bF_buf2), .C(_2581_), .Y(_2391_) );
	OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_25__28_), .Y(_2582_) );
	OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf3), .B(_2552__bF_buf1), .C(_2582_), .Y(_2392_) );
	OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_25__29_), .Y(_2583_) );
	OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf3), .B(_2552__bF_buf0), .C(_2583_), .Y(_2393_) );
	OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_25__30_), .Y(_2584_) );
	OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_2552__bF_buf4), .C(_2584_), .Y(_2394_) );
	OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_25__31_), .Y(_2585_) );
	OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf3), .B(_2552__bF_buf3), .C(_2585_), .Y(_2395_) );
	NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(biu_ins_7_), .Y(_2586_) );
	INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .Y(_2587_) );
	AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2587_), .Y(_2588_) );
	NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2480_), .C(_2588__bF_buf7), .Y(_2589_) );
	NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(biu_ins_7_), .C(_2469_), .Y(_2590_) );
	OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_26__0_), .Y(_2591_) );
	OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf2), .B(_2589__bF_buf4), .C(_2591_), .Y(_2396_) );
	OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_26__1_), .Y(_2592_) );
	OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf2), .B(_2589__bF_buf3), .C(_2592_), .Y(_2397_) );
	OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_26__2_), .Y(_2593_) );
	OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf2), .B(_2589__bF_buf2), .C(_2593_), .Y(_2398_) );
	OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_26__3_), .Y(_2594_) );
	OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf2), .B(_2589__bF_buf1), .C(_2594_), .Y(_2399_) );
	OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_26__4_), .Y(_2595_) );
	OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf2), .B(_2589__bF_buf0), .C(_2595_), .Y(_2400_) );
	OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_26__5_), .Y(_2596_) );
	OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf2), .B(_2589__bF_buf4), .C(_2596_), .Y(_2401_) );
	OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_26__6_), .Y(_2597_) );
	OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf2), .B(_2589__bF_buf3), .C(_2597_), .Y(_2402_) );
	OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_26__7_), .Y(_2598_) );
	OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf2), .B(_2589__bF_buf2), .C(_2598_), .Y(_2403_) );
	OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_26__8_), .Y(_2599_) );
	OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf2), .B(_2589__bF_buf1), .C(_2599_), .Y(_2404_) );
	OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_26__9_), .Y(_2600_) );
	OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf2), .B(_2589__bF_buf0), .C(_2600_), .Y(_2405_) );
	OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_26__10_), .Y(_2601_) );
	OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf2), .B(_2589__bF_buf4), .C(_2601_), .Y(_2406_) );
	OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_26__11_), .Y(_2602_) );
	OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf2), .B(_2589__bF_buf3), .C(_2602_), .Y(_2407_) );
	OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_26__12_), .Y(_2603_) );
	OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf2), .B(_2589__bF_buf2), .C(_2603_), .Y(_2408_) );
	OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_26__13_), .Y(_2604_) );
	OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf2), .B(_2589__bF_buf1), .C(_2604_), .Y(_2409_) );
	OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_26__14_), .Y(_2605_) );
	OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf2), .B(_2589__bF_buf0), .C(_2605_), .Y(_2410_) );
	OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_26__15_), .Y(_2606_) );
	OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf2), .B(_2589__bF_buf4), .C(_2606_), .Y(_2411_) );
	OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_26__16_), .Y(_2607_) );
	OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf2), .B(_2589__bF_buf3), .C(_2607_), .Y(_2412_) );
	OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_26__17_), .Y(_2608_) );
	OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf2), .B(_2589__bF_buf2), .C(_2608_), .Y(_2413_) );
	OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_26__18_), .Y(_2609_) );
	OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf2), .B(_2589__bF_buf1), .C(_2609_), .Y(_2414_) );
	OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_26__19_), .Y(_2610_) );
	OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf2), .B(_2589__bF_buf0), .C(_2610_), .Y(_2415_) );
	OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_26__20_), .Y(_2611_) );
	OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf2), .B(_2589__bF_buf4), .C(_2611_), .Y(_2416_) );
	OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_26__21_), .Y(_2612_) );
	OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf2), .B(_2589__bF_buf3), .C(_2612_), .Y(_2417_) );
	OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_26__22_), .Y(_2613_) );
	OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf2), .B(_2589__bF_buf2), .C(_2613_), .Y(_2418_) );
	OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_26__23_), .Y(_2614_) );
	OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf2), .B(_2589__bF_buf1), .C(_2614_), .Y(_2419_) );
	OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_26__24_), .Y(_2615_) );
	OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf2), .B(_2589__bF_buf0), .C(_2615_), .Y(_2420_) );
	OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_26__25_), .Y(_2616_) );
	OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf2), .B(_2589__bF_buf4), .C(_2616_), .Y(_2421_) );
	OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_26__26_), .Y(_2617_) );
	OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf2), .B(_2589__bF_buf3), .C(_2617_), .Y(_2422_) );
	OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_26__27_), .Y(_2618_) );
	OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf2), .B(_2589__bF_buf2), .C(_2618_), .Y(_2423_) );
	OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_26__28_), .Y(_2619_) );
	OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf2), .B(_2589__bF_buf1), .C(_2619_), .Y(_2424_) );
	OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_26__29_), .Y(_2620_) );
	OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf2), .B(_2589__bF_buf0), .C(_2620_), .Y(_2425_) );
	OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_26__30_), .Y(_2621_) );
	OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_2589__bF_buf4), .C(_2621_), .Y(_2426_) );
	OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_26__31_), .Y(_2622_) );
	OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf2), .B(_2589__bF_buf3), .C(_2622_), .Y(_2427_) );
	AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2461_), .Y(_2623_) );
	NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2480_), .C(_2623_), .Y(_2624_) );
	NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2469_), .Y(_2625_) );
	OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_27__0_), .Y(_2626_) );
	OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf1), .B(_2624__bF_buf4), .C(_2626_), .Y(_2428_) );
	OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_27__1_), .Y(_2627_) );
	OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf1), .B(_2624__bF_buf3), .C(_2627_), .Y(_2429_) );
	OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_27__2_), .Y(_2628_) );
	OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf1), .B(_2624__bF_buf2), .C(_2628_), .Y(_2430_) );
	OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_27__3_), .Y(_2629_) );
	OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf1), .B(_2624__bF_buf1), .C(_2629_), .Y(_2431_) );
	OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_27__4_), .Y(_2630_) );
	OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf1), .B(_2624__bF_buf0), .C(_2630_), .Y(_2432_) );
	OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_27__5_), .Y(_2631_) );
	OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf1), .B(_2624__bF_buf4), .C(_2631_), .Y(_2433_) );
	OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_27__6_), .Y(_2632_) );
	OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf1), .B(_2624__bF_buf3), .C(_2632_), .Y(_2434_) );
	OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_27__7_), .Y(_2633_) );
	OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf1), .B(_2624__bF_buf2), .C(_2633_), .Y(_2435_) );
	OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_27__8_), .Y(_2634_) );
	OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf1), .B(_2624__bF_buf1), .C(_2634_), .Y(_2436_) );
	OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_27__9_), .Y(_2635_) );
	OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf1), .B(_2624__bF_buf0), .C(_2635_), .Y(_2437_) );
	OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_27__10_), .Y(_2636_) );
	OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf1), .B(_2624__bF_buf4), .C(_2636_), .Y(_2438_) );
	OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_27__11_), .Y(_2637_) );
	OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf1), .B(_2624__bF_buf3), .C(_2637_), .Y(_2439_) );
	OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_27__12_), .Y(_2638_) );
	OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf1), .B(_2624__bF_buf2), .C(_2638_), .Y(_2440_) );
	OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_27__13_), .Y(_2639_) );
	OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf1), .B(_2624__bF_buf1), .C(_2639_), .Y(_2441_) );
	OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_27__14_), .Y(_2640_) );
	OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf1), .B(_2624__bF_buf0), .C(_2640_), .Y(_2442_) );
	OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_27__15_), .Y(_2641_) );
	OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf1), .B(_2624__bF_buf4), .C(_2641_), .Y(_2443_) );
	OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_27__16_), .Y(_2642_) );
	OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf1), .B(_2624__bF_buf3), .C(_2642_), .Y(_2444_) );
	OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_27__17_), .Y(_2643_) );
	OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf1), .B(_2624__bF_buf2), .C(_2643_), .Y(_2445_) );
	OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_27__18_), .Y(_2644_) );
	OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf1), .B(_2624__bF_buf1), .C(_2644_), .Y(_2446_) );
	OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_27__19_), .Y(_2645_) );
	OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf1), .B(_2624__bF_buf0), .C(_2645_), .Y(_2447_) );
	OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_27__20_), .Y(_2646_) );
	OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf1), .B(_2624__bF_buf4), .C(_2646_), .Y(_2448_) );
	OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_27__21_), .Y(_2647_) );
	OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf1), .B(_2624__bF_buf3), .C(_2647_), .Y(_2449_) );
	OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_27__22_), .Y(_2648_) );
	OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf1), .B(_2624__bF_buf2), .C(_2648_), .Y(_2450_) );
	OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_27__23_), .Y(_2649_) );
	OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf1), .B(_2624__bF_buf1), .C(_2649_), .Y(_2451_) );
	OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_27__24_), .Y(_2650_) );
	OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf1), .B(_2624__bF_buf0), .C(_2650_), .Y(_2452_) );
	OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_27__25_), .Y(_2651_) );
	OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf1), .B(_2624__bF_buf4), .C(_2651_), .Y(_2453_) );
	OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_27__26_), .Y(_2652_) );
	OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf1), .B(_2624__bF_buf3), .C(_2652_), .Y(_2454_) );
	OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_27__27_), .Y(_2653_) );
	OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf1), .B(_2624__bF_buf2), .C(_2653_), .Y(_2455_) );
	OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_27__28_), .Y(_2654_) );
	OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf1), .B(_2624__bF_buf1), .C(_2654_), .Y(_2456_) );
	OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_27__29_), .Y(_2655_) );
	OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf1), .B(_2624__bF_buf0), .C(_2655_), .Y(_2457_) );
	OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_27__30_), .Y(_2656_) );
	OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_2624__bF_buf4), .C(_2656_), .Y(_2458_) );
	OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_27__31_), .Y(_2657_) );
	OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf1), .B(_2624__bF_buf3), .C(_2657_), .Y(_2459_) );
	NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2480_), .C(_2588__bF_buf6), .Y(_2658_) );
	OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_30__0_), .Y(_2659_) );
	OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf0), .B(_2658__bF_buf4), .C(_2659_), .Y(_1468_) );
	OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_30__1_), .Y(_2660_) );
	OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf0), .B(_2658__bF_buf3), .C(_2660_), .Y(_1469_) );
	OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_30__2_), .Y(_2661_) );
	OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf0), .B(_2658__bF_buf2), .C(_2661_), .Y(_1470_) );
	OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_30__3_), .Y(_2662_) );
	OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf0), .B(_2658__bF_buf1), .C(_2662_), .Y(_1471_) );
	OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_30__4_), .Y(_2663_) );
	OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf0), .B(_2658__bF_buf0), .C(_2663_), .Y(_1472_) );
	OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_30__5_), .Y(_2664_) );
	OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf0), .B(_2658__bF_buf4), .C(_2664_), .Y(_1473_) );
	OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_30__6_), .Y(_2665_) );
	OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf0), .B(_2658__bF_buf3), .C(_2665_), .Y(_1474_) );
	OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_30__7_), .Y(_2666_) );
	OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf0), .B(_2658__bF_buf2), .C(_2666_), .Y(_1475_) );
	OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_30__8_), .Y(_2667_) );
	OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf0), .B(_2658__bF_buf1), .C(_2667_), .Y(_1476_) );
	OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_30__9_), .Y(_2668_) );
	OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf0), .B(_2658__bF_buf0), .C(_2668_), .Y(_1477_) );
	OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_30__10_), .Y(_2669_) );
	OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf0), .B(_2658__bF_buf4), .C(_2669_), .Y(_1478_) );
	OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_30__11_), .Y(_2670_) );
	OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf0), .B(_2658__bF_buf3), .C(_2670_), .Y(_1479_) );
	OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_30__12_), .Y(_2671_) );
	OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf0), .B(_2658__bF_buf2), .C(_2671_), .Y(_1480_) );
	OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_30__13_), .Y(_2672_) );
	OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf0), .B(_2658__bF_buf1), .C(_2672_), .Y(_1481_) );
	OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_30__14_), .Y(_2673_) );
	OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf0), .B(_2658__bF_buf0), .C(_2673_), .Y(_1482_) );
	OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_30__15_), .Y(_2674_) );
	OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf0), .B(_2658__bF_buf4), .C(_2674_), .Y(_1483_) );
	OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_30__16_), .Y(_2675_) );
	OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf0), .B(_2658__bF_buf3), .C(_2675_), .Y(_1484_) );
	OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_30__17_), .Y(_2676_) );
	OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf0), .B(_2658__bF_buf2), .C(_2676_), .Y(_1485_) );
	OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_30__18_), .Y(_2677_) );
	OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf0), .B(_2658__bF_buf1), .C(_2677_), .Y(_1486_) );
	OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_30__19_), .Y(_2678_) );
	OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf0), .B(_2658__bF_buf0), .C(_2678_), .Y(_1487_) );
	OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_30__20_), .Y(_2679_) );
	OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf0), .B(_2658__bF_buf4), .C(_2679_), .Y(_1488_) );
	OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_30__21_), .Y(_2680_) );
	OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf0), .B(_2658__bF_buf3), .C(_2680_), .Y(_1489_) );
	OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_30__22_), .Y(_2681_) );
	OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf0), .B(_2658__bF_buf2), .C(_2681_), .Y(_1490_) );
	OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_30__23_), .Y(_2682_) );
	OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf0), .B(_2658__bF_buf1), .C(_2682_), .Y(_1491_) );
	OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_30__24_), .Y(_2683_) );
	OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf0), .B(_2658__bF_buf0), .C(_2683_), .Y(_1492_) );
	OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_30__25_), .Y(_2684_) );
	OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf0), .B(_2658__bF_buf4), .C(_2684_), .Y(_1493_) );
	OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_30__26_), .Y(_2685_) );
	OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf0), .B(_2658__bF_buf3), .C(_2685_), .Y(_1494_) );
	OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_30__27_), .Y(_2686_) );
	OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf0), .B(_2658__bF_buf2), .C(_2686_), .Y(_1495_) );
	OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_30__28_), .Y(_2687_) );
	OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf0), .B(_2658__bF_buf1), .C(_2687_), .Y(_1496_) );
	OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_30__29_), .Y(_2688_) );
	OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf0), .B(_2658__bF_buf0), .C(_2688_), .Y(_1497_) );
	OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_30__30_), .Y(_2689_) );
	OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_2658__bF_buf4), .C(_2689_), .Y(_1498_) );
	OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_30__31_), .Y(_2690_) );
	OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf0), .B(_2658__bF_buf3), .C(_2690_), .Y(_1499_) );
	INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .Y(_2691_) );
	NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_7_), .B(_2691_), .Y(_2692_) );
	INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(_2692_), .Y(_2693_) );
	AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2693_), .Y(_2694_) );
	NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2480_), .C(_2694__bF_buf7), .Y(_2695_) );
	NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(biu_ins_7_), .C(_2469_), .Y(_2696_) );
	OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_28__0_), .Y(_2697_) );
	OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf4), .B(_2695__bF_buf4), .C(_2697_), .Y(_1500_) );
	OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_28__1_), .Y(_2698_) );
	OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf4), .B(_2695__bF_buf3), .C(_2698_), .Y(_1501_) );
	OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_28__2_), .Y(_2699_) );
	OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf4), .B(_2695__bF_buf2), .C(_2699_), .Y(_1502_) );
	OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_28__3_), .Y(_2700_) );
	OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf4), .B(_2695__bF_buf1), .C(_2700_), .Y(_1503_) );
	OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_28__4_), .Y(_2701_) );
	OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf4), .B(_2695__bF_buf0), .C(_2701_), .Y(_1504_) );
	OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_28__5_), .Y(_2702_) );
	OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf4), .B(_2695__bF_buf4), .C(_2702_), .Y(_1505_) );
	OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_28__6_), .Y(_2703_) );
	OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf4), .B(_2695__bF_buf3), .C(_2703_), .Y(_1506_) );
	OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_28__7_), .Y(_2704_) );
	OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf4), .B(_2695__bF_buf2), .C(_2704_), .Y(_1507_) );
	OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_28__8_), .Y(_2705_) );
	OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf4), .B(_2695__bF_buf1), .C(_2705_), .Y(_1508_) );
	OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_28__9_), .Y(_2706_) );
	OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf4), .B(_2695__bF_buf0), .C(_2706_), .Y(_1509_) );
	OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_28__10_), .Y(_2707_) );
	OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf4), .B(_2695__bF_buf4), .C(_2707_), .Y(_1510_) );
	OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_28__11_), .Y(_2708_) );
	OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf4), .B(_2695__bF_buf3), .C(_2708_), .Y(_1511_) );
	OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_28__12_), .Y(_2709_) );
	OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf4), .B(_2695__bF_buf2), .C(_2709_), .Y(_1512_) );
	OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_28__13_), .Y(_2710_) );
	OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf4), .B(_2695__bF_buf1), .C(_2710_), .Y(_1513_) );
	OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_28__14_), .Y(_2711_) );
	OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf4), .B(_2695__bF_buf0), .C(_2711_), .Y(_1514_) );
	OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_28__15_), .Y(_2712_) );
	OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf4), .B(_2695__bF_buf4), .C(_2712_), .Y(_1515_) );
	OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_28__16_), .Y(_2713_) );
	OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf4), .B(_2695__bF_buf3), .C(_2713_), .Y(_1516_) );
	OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_28__17_), .Y(_2714_) );
	OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf4), .B(_2695__bF_buf2), .C(_2714_), .Y(_1517_) );
	OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_28__18_), .Y(_2715_) );
	OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf4), .B(_2695__bF_buf1), .C(_2715_), .Y(_1518_) );
	OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_28__19_), .Y(_2716_) );
	OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf4), .B(_2695__bF_buf0), .C(_2716_), .Y(_1519_) );
	OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_28__20_), .Y(_2717_) );
	OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf4), .B(_2695__bF_buf4), .C(_2717_), .Y(_1520_) );
	OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_28__21_), .Y(_2718_) );
	OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf4), .B(_2695__bF_buf3), .C(_2718_), .Y(_1521_) );
	OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_28__22_), .Y(_2719_) );
	OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf4), .B(_2695__bF_buf2), .C(_2719_), .Y(_1522_) );
	OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_2487__bF_buf2), .C(csr_gpr_iu_gpr_28__23_), .Y(_2720_) );
	OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf4), .B(_2695__bF_buf1), .C(_2720_), .Y(_1523_) );
	OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_2487__bF_buf1), .C(csr_gpr_iu_gpr_28__24_), .Y(_2721_) );
	OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf4), .B(_2695__bF_buf0), .C(_2721_), .Y(_1524_) );
	OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_2487__bF_buf0), .C(csr_gpr_iu_gpr_28__25_), .Y(_2722_) );
	OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf4), .B(_2695__bF_buf4), .C(_2722_), .Y(_1525_) );
	OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_2487__bF_buf8), .C(csr_gpr_iu_gpr_28__26_), .Y(_2723_) );
	OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf4), .B(_2695__bF_buf3), .C(_2723_), .Y(_1526_) );
	OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_2487__bF_buf7), .C(csr_gpr_iu_gpr_28__27_), .Y(_2724_) );
	OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf4), .B(_2695__bF_buf2), .C(_2724_), .Y(_1527_) );
	OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_2487__bF_buf6), .C(csr_gpr_iu_gpr_28__28_), .Y(_2725_) );
	OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf4), .B(_2695__bF_buf1), .C(_2725_), .Y(_1528_) );
	OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_2487__bF_buf5), .C(csr_gpr_iu_gpr_28__29_), .Y(_2726_) );
	OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf4), .B(_2695__bF_buf0), .C(_2726_), .Y(_1529_) );
	OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_2487__bF_buf4), .C(csr_gpr_iu_gpr_28__30_), .Y(_2727_) );
	OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_2695__bF_buf4), .C(_2727_), .Y(_1530_) );
	OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_2487__bF_buf3), .C(csr_gpr_iu_gpr_28__31_), .Y(_2728_) );
	OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf4), .B(_2695__bF_buf3), .C(_2728_), .Y(_1531_) );
	INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__0_), .Y(_2729_) );
	NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2479_), .C(_2482_), .Y(_2730_) );
	NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2696__bF_buf6), .Y(_2731_) );
	INVX8 INVX8_45 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .Y(_2732_) );
	NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2732__bF_buf8), .C(_2694__bF_buf6), .Y(_2733_) );
	OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_2729_), .B(_2731__bF_buf4), .C(_2733_), .Y(_1532_) );
	INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__1_), .Y(_2734_) );
	NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2732__bF_buf7), .C(_2694__bF_buf5), .Y(_2735_) );
	OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_2731__bF_buf3), .C(_2735_), .Y(_1533_) );
	INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__2_), .Y(_2736_) );
	NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2732__bF_buf6), .C(_2694__bF_buf4), .Y(_2737_) );
	OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(_2731__bF_buf2), .C(_2737_), .Y(_1534_) );
	INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__3_), .Y(_2738_) );
	NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2732__bF_buf5), .C(_2694__bF_buf3), .Y(_2739_) );
	OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2731__bF_buf1), .C(_2739_), .Y(_1535_) );
	INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__4_), .Y(_2740_) );
	NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2732__bF_buf4), .C(_2694__bF_buf2), .Y(_2741_) );
	OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .B(_2731__bF_buf0), .C(_2741_), .Y(_1536_) );
	INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__5_), .Y(_2742_) );
	NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2732__bF_buf3), .C(_2694__bF_buf1), .Y(_2743_) );
	OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2731__bF_buf4), .C(_2743_), .Y(_1537_) );
	INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__6_), .Y(_2744_) );
	NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2732__bF_buf2), .C(_2694__bF_buf0), .Y(_2745_) );
	OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_2744_), .B(_2731__bF_buf3), .C(_2745_), .Y(_1538_) );
	INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__7_), .Y(_2746_) );
	NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2732__bF_buf1), .C(_2694__bF_buf7), .Y(_2747_) );
	OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_2746_), .B(_2731__bF_buf2), .C(_2747_), .Y(_1539_) );
	INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__8_), .Y(_2748_) );
	NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2732__bF_buf0), .C(_2694__bF_buf6), .Y(_2749_) );
	OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2731__bF_buf1), .C(_2749_), .Y(_1540_) );
	INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__9_), .Y(_2750_) );
	NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2732__bF_buf8), .C(_2694__bF_buf5), .Y(_2751_) );
	OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_2731__bF_buf0), .C(_2751_), .Y(_1541_) );
	INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__10_), .Y(_2752_) );
	NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2732__bF_buf7), .C(_2694__bF_buf4), .Y(_2753_) );
	OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_2752_), .B(_2731__bF_buf4), .C(_2753_), .Y(_1542_) );
	INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__11_), .Y(_2754_) );
	NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2732__bF_buf6), .C(_2694__bF_buf3), .Y(_2755_) );
	OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2731__bF_buf3), .C(_2755_), .Y(_1543_) );
	INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__12_), .Y(_2756_) );
	NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2732__bF_buf5), .C(_2694__bF_buf2), .Y(_2757_) );
	OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_2731__bF_buf2), .C(_2757_), .Y(_1544_) );
	INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__13_), .Y(_2758_) );
	NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2732__bF_buf4), .C(_2694__bF_buf1), .Y(_2759_) );
	OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_2758_), .B(_2731__bF_buf1), .C(_2759_), .Y(_1545_) );
	INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__14_), .Y(_2760_) );
	NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2732__bF_buf3), .C(_2694__bF_buf0), .Y(_2761_) );
	OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2731__bF_buf0), .C(_2761_), .Y(_1546_) );
	INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__15_), .Y(_2762_) );
	NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2732__bF_buf2), .C(_2694__bF_buf7), .Y(_2763_) );
	OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_2731__bF_buf4), .C(_2763_), .Y(_1547_) );
	INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__16_), .Y(_2764_) );
	NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2732__bF_buf1), .C(_2694__bF_buf6), .Y(_2765_) );
	OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_2764_), .B(_2731__bF_buf3), .C(_2765_), .Y(_1548_) );
	INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__17_), .Y(_2766_) );
	NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2732__bF_buf0), .C(_2694__bF_buf5), .Y(_2767_) );
	OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2731__bF_buf2), .C(_2767_), .Y(_1549_) );
	INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__18_), .Y(_2768_) );
	NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2732__bF_buf8), .C(_2694__bF_buf4), .Y(_2769_) );
	OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_2731__bF_buf1), .C(_2769_), .Y(_1550_) );
	INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__19_), .Y(_2770_) );
	NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2732__bF_buf7), .C(_2694__bF_buf3), .Y(_2771_) );
	OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_2770_), .B(_2731__bF_buf0), .C(_2771_), .Y(_1551_) );
	INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__20_), .Y(_2772_) );
	NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2732__bF_buf6), .C(_2694__bF_buf2), .Y(_2773_) );
	OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_2731__bF_buf4), .C(_2773_), .Y(_1552_) );
	INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__21_), .Y(_2774_) );
	NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2732__bF_buf5), .C(_2694__bF_buf1), .Y(_2775_) );
	OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .B(_2731__bF_buf3), .C(_2775_), .Y(_1553_) );
	INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__22_), .Y(_2776_) );
	NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2732__bF_buf4), .C(_2694__bF_buf0), .Y(_2777_) );
	OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2731__bF_buf2), .C(_2777_), .Y(_1554_) );
	INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__23_), .Y(_2778_) );
	NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2732__bF_buf3), .C(_2694__bF_buf7), .Y(_2779_) );
	OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_2778_), .B(_2731__bF_buf1), .C(_2779_), .Y(_1555_) );
	INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__24_), .Y(_2780_) );
	NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2732__bF_buf2), .C(_2694__bF_buf6), .Y(_2781_) );
	OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_2731__bF_buf0), .C(_2781_), .Y(_1556_) );
	INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__25_), .Y(_2782_) );
	NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2732__bF_buf1), .C(_2694__bF_buf5), .Y(_2783_) );
	OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_2782_), .B(_2731__bF_buf4), .C(_2783_), .Y(_1557_) );
	INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__26_), .Y(_2784_) );
	NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2732__bF_buf0), .C(_2694__bF_buf4), .Y(_2785_) );
	OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_2784_), .B(_2731__bF_buf3), .C(_2785_), .Y(_1558_) );
	INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__27_), .Y(_2786_) );
	NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2732__bF_buf8), .C(_2694__bF_buf3), .Y(_2787_) );
	OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2731__bF_buf2), .C(_2787_), .Y(_1559_) );
	INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__28_), .Y(_2788_) );
	NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2732__bF_buf7), .C(_2694__bF_buf2), .Y(_2789_) );
	OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2731__bF_buf1), .C(_2789_), .Y(_1560_) );
	INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__29_), .Y(_2790_) );
	NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2732__bF_buf6), .C(_2694__bF_buf1), .Y(_2791_) );
	OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2731__bF_buf0), .C(_2791_), .Y(_1561_) );
	INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__30_), .Y(_2792_) );
	NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2732__bF_buf5), .C(_2694__bF_buf0), .Y(_2793_) );
	OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_2792_), .B(_2731__bF_buf4), .C(_2793_), .Y(_1562_) );
	INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_20__31_), .Y(_2794_) );
	NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2732__bF_buf4), .C(_2694__bF_buf7), .Y(_2795_) );
	OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .B(_2731__bF_buf3), .C(_2795_), .Y(_1563_) );
	INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__0_), .Y(_2796_) );
	NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2484__bF_buf0), .Y(_2797_) );
	NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2732__bF_buf3), .C(_2473__bF_buf5), .Y(_2798_) );
	OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_2796_), .B(_2797__bF_buf4), .C(_2798_), .Y(_1564_) );
	INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__1_), .Y(_2799_) );
	NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2732__bF_buf2), .C(_2473__bF_buf4), .Y(_2800_) );
	OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_2797__bF_buf3), .C(_2800_), .Y(_1565_) );
	INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__2_), .Y(_2801_) );
	NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2732__bF_buf1), .C(_2473__bF_buf3), .Y(_2802_) );
	OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_2801_), .B(_2797__bF_buf2), .C(_2802_), .Y(_1566_) );
	INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__3_), .Y(_2803_) );
	NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2732__bF_buf0), .C(_2473__bF_buf2), .Y(_2804_) );
	OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_2797__bF_buf1), .C(_2804_), .Y(_1567_) );
	INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__4_), .Y(_2805_) );
	NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2732__bF_buf8), .C(_2473__bF_buf1), .Y(_2806_) );
	OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_2797__bF_buf0), .C(_2806_), .Y(_1568_) );
	INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__5_), .Y(_2807_) );
	NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2732__bF_buf7), .C(_2473__bF_buf0), .Y(_2808_) );
	OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .B(_2797__bF_buf4), .C(_2808_), .Y(_1569_) );
	INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__6_), .Y(_2809_) );
	NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2732__bF_buf6), .C(_2473__bF_buf7), .Y(_2810_) );
	OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_2809_), .B(_2797__bF_buf3), .C(_2810_), .Y(_1570_) );
	INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__7_), .Y(_2811_) );
	NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2732__bF_buf5), .C(_2473__bF_buf6), .Y(_2812_) );
	OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_2811_), .B(_2797__bF_buf2), .C(_2812_), .Y(_1571_) );
	INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__8_), .Y(_2813_) );
	NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2732__bF_buf4), .C(_2473__bF_buf5), .Y(_2814_) );
	OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_2797__bF_buf1), .C(_2814_), .Y(_1572_) );
	INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__9_), .Y(_2815_) );
	NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2732__bF_buf3), .C(_2473__bF_buf4), .Y(_2816_) );
	OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_2797__bF_buf0), .C(_2816_), .Y(_1573_) );
	INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__10_), .Y(_2817_) );
	NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2732__bF_buf2), .C(_2473__bF_buf3), .Y(_2818_) );
	OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(_2797__bF_buf4), .C(_2818_), .Y(_1574_) );
	INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__11_), .Y(_2819_) );
	NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2732__bF_buf1), .C(_2473__bF_buf2), .Y(_2820_) );
	OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .B(_2797__bF_buf3), .C(_2820_), .Y(_1575_) );
	INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__12_), .Y(_2821_) );
	NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2732__bF_buf0), .C(_2473__bF_buf1), .Y(_2822_) );
	OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_2797__bF_buf2), .C(_2822_), .Y(_1576_) );
	INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__13_), .Y(_2823_) );
	NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2732__bF_buf8), .C(_2473__bF_buf0), .Y(_2824_) );
	OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_2797__bF_buf1), .C(_2824_), .Y(_1577_) );
	INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__14_), .Y(_2825_) );
	NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2732__bF_buf7), .C(_2473__bF_buf7), .Y(_2826_) );
	OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_2797__bF_buf0), .C(_2826_), .Y(_1578_) );
	INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__15_), .Y(_2827_) );
	NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2732__bF_buf6), .C(_2473__bF_buf6), .Y(_2828_) );
	OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_2797__bF_buf4), .C(_2828_), .Y(_1579_) );
	INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__16_), .Y(_2829_) );
	NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2732__bF_buf5), .C(_2473__bF_buf5), .Y(_2830_) );
	OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_2829_), .B(_2797__bF_buf3), .C(_2830_), .Y(_1580_) );
	INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__17_), .Y(_2831_) );
	NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2732__bF_buf4), .C(_2473__bF_buf4), .Y(_2832_) );
	OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_2797__bF_buf2), .C(_2832_), .Y(_1581_) );
	INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__18_), .Y(_2833_) );
	NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2732__bF_buf3), .C(_2473__bF_buf3), .Y(_2834_) );
	OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .B(_2797__bF_buf1), .C(_2834_), .Y(_1582_) );
	INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__19_), .Y(_2835_) );
	NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2732__bF_buf2), .C(_2473__bF_buf2), .Y(_2836_) );
	OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .B(_2797__bF_buf0), .C(_2836_), .Y(_1583_) );
	INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__20_), .Y(_2837_) );
	NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2732__bF_buf1), .C(_2473__bF_buf1), .Y(_2838_) );
	OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .B(_2797__bF_buf4), .C(_2838_), .Y(_1584_) );
	INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__21_), .Y(_2839_) );
	NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2732__bF_buf0), .C(_2473__bF_buf0), .Y(_2840_) );
	OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_2797__bF_buf3), .C(_2840_), .Y(_1585_) );
	INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__22_), .Y(_2841_) );
	NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2732__bF_buf8), .C(_2473__bF_buf7), .Y(_2842_) );
	OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_2841_), .B(_2797__bF_buf2), .C(_2842_), .Y(_1586_) );
	INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__23_), .Y(_2843_) );
	NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2732__bF_buf7), .C(_2473__bF_buf6), .Y(_2844_) );
	OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_2843_), .B(_2797__bF_buf1), .C(_2844_), .Y(_1587_) );
	INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__24_), .Y(_2845_) );
	NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2732__bF_buf6), .C(_2473__bF_buf5), .Y(_2846_) );
	OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_2845_), .B(_2797__bF_buf0), .C(_2846_), .Y(_1588_) );
	INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__25_), .Y(_2847_) );
	NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2732__bF_buf5), .C(_2473__bF_buf4), .Y(_2848_) );
	OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_2797__bF_buf4), .C(_2848_), .Y(_1589_) );
	INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__26_), .Y(_2849_) );
	NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2732__bF_buf4), .C(_2473__bF_buf3), .Y(_2850_) );
	OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_2797__bF_buf3), .C(_2850_), .Y(_1590_) );
	INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__27_), .Y(_2851_) );
	NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2732__bF_buf3), .C(_2473__bF_buf2), .Y(_2852_) );
	OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_2851_), .B(_2797__bF_buf2), .C(_2852_), .Y(_1591_) );
	INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__28_), .Y(_2853_) );
	NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2732__bF_buf2), .C(_2473__bF_buf1), .Y(_2854_) );
	OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2797__bF_buf1), .C(_2854_), .Y(_1592_) );
	INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__29_), .Y(_2855_) );
	NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2732__bF_buf1), .C(_2473__bF_buf0), .Y(_2856_) );
	OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2797__bF_buf0), .C(_2856_), .Y(_1593_) );
	INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__30_), .Y(_2857_) );
	NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2732__bF_buf0), .C(_2473__bF_buf7), .Y(_2858_) );
	OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_2797__bF_buf4), .C(_2858_), .Y(_1594_) );
	INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_21__31_), .Y(_2859_) );
	NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2732__bF_buf8), .C(_2473__bF_buf6), .Y(_2860_) );
	OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_2797__bF_buf3), .C(_2860_), .Y(_1595_) );
	INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__0_), .Y(_2861_) );
	NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2590__bF_buf0), .Y(_2862_) );
	NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2732__bF_buf7), .C(_2588__bF_buf5), .Y(_2863_) );
	OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_2862__bF_buf4), .C(_2863_), .Y(_1596_) );
	INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__1_), .Y(_2864_) );
	NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2732__bF_buf6), .C(_2588__bF_buf4), .Y(_2865_) );
	OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_2862__bF_buf3), .C(_2865_), .Y(_1597_) );
	INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__2_), .Y(_2866_) );
	NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2732__bF_buf5), .C(_2588__bF_buf3), .Y(_2867_) );
	OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_2862__bF_buf2), .C(_2867_), .Y(_1598_) );
	INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__3_), .Y(_2868_) );
	NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2732__bF_buf4), .C(_2588__bF_buf2), .Y(_2869_) );
	OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(_2862__bF_buf1), .C(_2869_), .Y(_1599_) );
	INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__4_), .Y(_2870_) );
	NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2732__bF_buf3), .C(_2588__bF_buf1), .Y(_2871_) );
	OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_2862__bF_buf0), .C(_2871_), .Y(_1600_) );
	INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__5_), .Y(_2872_) );
	NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2732__bF_buf2), .C(_2588__bF_buf0), .Y(_2873_) );
	OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2862__bF_buf4), .C(_2873_), .Y(_1601_) );
	INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__6_), .Y(_2874_) );
	NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2732__bF_buf1), .C(_2588__bF_buf7), .Y(_2875_) );
	OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .B(_2862__bF_buf3), .C(_2875_), .Y(_1602_) );
	INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__7_), .Y(_2876_) );
	NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2732__bF_buf0), .C(_2588__bF_buf6), .Y(_2877_) );
	OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_2862__bF_buf2), .C(_2877_), .Y(_1603_) );
	INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__8_), .Y(_2878_) );
	NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2732__bF_buf8), .C(_2588__bF_buf5), .Y(_2879_) );
	OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_2862__bF_buf1), .C(_2879_), .Y(_1604_) );
	INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__9_), .Y(_2880_) );
	NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2732__bF_buf7), .C(_2588__bF_buf4), .Y(_2881_) );
	OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_2862__bF_buf0), .C(_2881_), .Y(_1605_) );
	INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__10_), .Y(_2882_) );
	NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2732__bF_buf6), .C(_2588__bF_buf3), .Y(_2883_) );
	OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_2862__bF_buf4), .C(_2883_), .Y(_1606_) );
	INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__11_), .Y(_2884_) );
	NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2732__bF_buf5), .C(_2588__bF_buf2), .Y(_2885_) );
	OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_2862__bF_buf3), .C(_2885_), .Y(_1607_) );
	INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__12_), .Y(_2886_) );
	NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2732__bF_buf4), .C(_2588__bF_buf1), .Y(_2887_) );
	OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .B(_2862__bF_buf2), .C(_2887_), .Y(_1608_) );
	INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__13_), .Y(_2888_) );
	NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2732__bF_buf3), .C(_2588__bF_buf0), .Y(_2889_) );
	OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_2862__bF_buf1), .C(_2889_), .Y(_1609_) );
	INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__14_), .Y(_2890_) );
	NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2732__bF_buf2), .C(_2588__bF_buf7), .Y(_2891_) );
	OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_2862__bF_buf0), .C(_2891_), .Y(_1610_) );
	INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__15_), .Y(_2892_) );
	NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2732__bF_buf1), .C(_2588__bF_buf6), .Y(_2893_) );
	OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_2892_), .B(_2862__bF_buf4), .C(_2893_), .Y(_1611_) );
	INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__16_), .Y(_2894_) );
	NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2732__bF_buf0), .C(_2588__bF_buf5), .Y(_2895_) );
	OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_2862__bF_buf3), .C(_2895_), .Y(_1612_) );
	INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__17_), .Y(_2896_) );
	NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2732__bF_buf8), .C(_2588__bF_buf4), .Y(_2897_) );
	OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_2862__bF_buf2), .C(_2897_), .Y(_1613_) );
	INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__18_), .Y(_2898_) );
	NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2732__bF_buf7), .C(_2588__bF_buf3), .Y(_2899_) );
	OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_2862__bF_buf1), .C(_2899_), .Y(_1614_) );
	INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__19_), .Y(_2900_) );
	NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2732__bF_buf6), .C(_2588__bF_buf2), .Y(_2901_) );
	OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_2862__bF_buf0), .C(_2901_), .Y(_1615_) );
	INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__20_), .Y(_2902_) );
	NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2732__bF_buf5), .C(_2588__bF_buf1), .Y(_2903_) );
	OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_2862__bF_buf4), .C(_2903_), .Y(_1616_) );
	INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__21_), .Y(_2904_) );
	NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2732__bF_buf4), .C(_2588__bF_buf0), .Y(_2905_) );
	OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(_2862__bF_buf3), .C(_2905_), .Y(_1617_) );
	INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__22_), .Y(_2906_) );
	NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2732__bF_buf3), .C(_2588__bF_buf7), .Y(_2907_) );
	OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .B(_2862__bF_buf2), .C(_2907_), .Y(_1618_) );
	INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__23_), .Y(_2908_) );
	NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2732__bF_buf2), .C(_2588__bF_buf6), .Y(_2909_) );
	OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_2862__bF_buf1), .C(_2909_), .Y(_1619_) );
	INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__24_), .Y(_2910_) );
	NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2732__bF_buf1), .C(_2588__bF_buf5), .Y(_2911_) );
	OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_2910_), .B(_2862__bF_buf0), .C(_2911_), .Y(_1620_) );
	INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__25_), .Y(_2912_) );
	NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2732__bF_buf0), .C(_2588__bF_buf4), .Y(_2913_) );
	OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_2862__bF_buf4), .C(_2913_), .Y(_1621_) );
	INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__26_), .Y(_2914_) );
	NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2732__bF_buf8), .C(_2588__bF_buf3), .Y(_2915_) );
	OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_2862__bF_buf3), .C(_2915_), .Y(_1622_) );
	INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__27_), .Y(_2916_) );
	NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2732__bF_buf7), .C(_2588__bF_buf2), .Y(_2917_) );
	OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .B(_2862__bF_buf2), .C(_2917_), .Y(_1623_) );
	INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__28_), .Y(_2918_) );
	NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2732__bF_buf6), .C(_2588__bF_buf1), .Y(_2919_) );
	OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .B(_2862__bF_buf1), .C(_2919_), .Y(_1624_) );
	INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__29_), .Y(_2920_) );
	NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2732__bF_buf5), .C(_2588__bF_buf0), .Y(_2921_) );
	OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2862__bF_buf0), .C(_2921_), .Y(_1625_) );
	INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__30_), .Y(_2922_) );
	NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2732__bF_buf4), .C(_2588__bF_buf7), .Y(_2923_) );
	OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_2862__bF_buf4), .C(_2923_), .Y(_1626_) );
	INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_22__31_), .Y(_2924_) );
	NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2732__bF_buf3), .C(_2588__bF_buf6), .Y(_2925_) );
	OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2862__bF_buf3), .C(_2925_), .Y(_1627_) );
	NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2732__bF_buf2), .B(_2623_), .Y(_2926_) );
	OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf12), .C(csr_gpr_iu_gpr_23__0_), .Y(_2927_) );
	OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf3), .B(_2926__bF_buf4), .C(_2927_), .Y(_1628_) );
	OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf11), .C(csr_gpr_iu_gpr_23__1_), .Y(_2928_) );
	OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf3), .B(_2926__bF_buf3), .C(_2928_), .Y(_1629_) );
	OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2625__bF_buf10), .C(csr_gpr_iu_gpr_23__2_), .Y(_2929_) );
	OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf3), .B(_2926__bF_buf2), .C(_2929_), .Y(_1630_) );
	OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .B(_2625__bF_buf9), .C(csr_gpr_iu_gpr_23__3_), .Y(_2930_) );
	OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf3), .B(_2926__bF_buf1), .C(_2930_), .Y(_1631_) );
	OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2625__bF_buf8), .C(csr_gpr_iu_gpr_23__4_), .Y(_2931_) );
	OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf3), .B(_2926__bF_buf0), .C(_2931_), .Y(_1632_) );
	OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2625__bF_buf7), .C(csr_gpr_iu_gpr_23__5_), .Y(_2932_) );
	OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf3), .B(_2926__bF_buf4), .C(_2932_), .Y(_1633_) );
	OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf6), .C(csr_gpr_iu_gpr_23__6_), .Y(_2933_) );
	OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf3), .B(_2926__bF_buf3), .C(_2933_), .Y(_1634_) );
	OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf5), .C(csr_gpr_iu_gpr_23__7_), .Y(_2934_) );
	OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf3), .B(_2926__bF_buf2), .C(_2934_), .Y(_1635_) );
	OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2625__bF_buf4), .C(csr_gpr_iu_gpr_23__8_), .Y(_2935_) );
	OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf3), .B(_2926__bF_buf1), .C(_2935_), .Y(_1636_) );
	OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .B(_2625__bF_buf3), .C(csr_gpr_iu_gpr_23__9_), .Y(_2936_) );
	OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf3), .B(_2926__bF_buf0), .C(_2936_), .Y(_1637_) );
	OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2625__bF_buf2), .C(csr_gpr_iu_gpr_23__10_), .Y(_2937_) );
	OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf3), .B(_2926__bF_buf4), .C(_2937_), .Y(_1638_) );
	OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2625__bF_buf1), .C(csr_gpr_iu_gpr_23__11_), .Y(_2938_) );
	OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf3), .B(_2926__bF_buf3), .C(_2938_), .Y(_1639_) );
	OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf0), .C(csr_gpr_iu_gpr_23__12_), .Y(_2939_) );
	OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf3), .B(_2926__bF_buf2), .C(_2939_), .Y(_1640_) );
	OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf14), .C(csr_gpr_iu_gpr_23__13_), .Y(_2940_) );
	OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf3), .B(_2926__bF_buf1), .C(_2940_), .Y(_1641_) );
	OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2625__bF_buf13), .C(csr_gpr_iu_gpr_23__14_), .Y(_2941_) );
	OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf3), .B(_2926__bF_buf0), .C(_2941_), .Y(_1642_) );
	OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .B(_2625__bF_buf12), .C(csr_gpr_iu_gpr_23__15_), .Y(_2942_) );
	OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf3), .B(_2926__bF_buf4), .C(_2942_), .Y(_1643_) );
	OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2625__bF_buf11), .C(csr_gpr_iu_gpr_23__16_), .Y(_2943_) );
	OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf3), .B(_2926__bF_buf3), .C(_2943_), .Y(_1644_) );
	OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2625__bF_buf10), .C(csr_gpr_iu_gpr_23__17_), .Y(_2944_) );
	OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf3), .B(_2926__bF_buf2), .C(_2944_), .Y(_1645_) );
	OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf9), .C(csr_gpr_iu_gpr_23__18_), .Y(_2945_) );
	OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf3), .B(_2926__bF_buf1), .C(_2945_), .Y(_1646_) );
	OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf8), .C(csr_gpr_iu_gpr_23__19_), .Y(_2946_) );
	OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf3), .B(_2926__bF_buf0), .C(_2946_), .Y(_1647_) );
	OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2625__bF_buf7), .C(csr_gpr_iu_gpr_23__20_), .Y(_2947_) );
	OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf3), .B(_2926__bF_buf4), .C(_2947_), .Y(_1648_) );
	OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .B(_2625__bF_buf6), .C(csr_gpr_iu_gpr_23__21_), .Y(_2948_) );
	OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf3), .B(_2926__bF_buf3), .C(_2948_), .Y(_1649_) );
	OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2625__bF_buf5), .C(csr_gpr_iu_gpr_23__22_), .Y(_2949_) );
	OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf3), .B(_2926__bF_buf2), .C(_2949_), .Y(_1650_) );
	OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2625__bF_buf4), .C(csr_gpr_iu_gpr_23__23_), .Y(_2950_) );
	OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf3), .B(_2926__bF_buf1), .C(_2950_), .Y(_1651_) );
	OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf3), .C(csr_gpr_iu_gpr_23__24_), .Y(_2951_) );
	OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf3), .B(_2926__bF_buf0), .C(_2951_), .Y(_1652_) );
	OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf2), .C(csr_gpr_iu_gpr_23__25_), .Y(_2952_) );
	OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf3), .B(_2926__bF_buf4), .C(_2952_), .Y(_1653_) );
	OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf5), .B(_2625__bF_buf1), .C(csr_gpr_iu_gpr_23__26_), .Y(_2953_) );
	OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf3), .B(_2926__bF_buf3), .C(_2953_), .Y(_1654_) );
	OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf4), .B(_2625__bF_buf0), .C(csr_gpr_iu_gpr_23__27_), .Y(_2954_) );
	OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf3), .B(_2926__bF_buf2), .C(_2954_), .Y(_1655_) );
	OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf3), .B(_2625__bF_buf14), .C(csr_gpr_iu_gpr_23__28_), .Y(_2955_) );
	OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf3), .B(_2926__bF_buf1), .C(_2955_), .Y(_1656_) );
	OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf2), .B(_2625__bF_buf13), .C(csr_gpr_iu_gpr_23__29_), .Y(_2956_) );
	OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf3), .B(_2926__bF_buf0), .C(_2956_), .Y(_1657_) );
	OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf1), .B(_2625__bF_buf12), .C(csr_gpr_iu_gpr_23__30_), .Y(_2957_) );
	OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_2926__bF_buf4), .C(_2957_), .Y(_1658_) );
	OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_2730__bF_buf0), .B(_2625__bF_buf11), .C(csr_gpr_iu_gpr_23__31_), .Y(_2958_) );
	OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf3), .B(_2926__bF_buf3), .C(_2958_), .Y(_1659_) );
	NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2480_), .C(_2694__bF_buf6), .Y(_2959_) );
	OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_24__0_), .Y(_2960_) );
	OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf2), .B(_2959__bF_buf4), .C(_2960_), .Y(_1660_) );
	OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_24__1_), .Y(_2961_) );
	OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf2), .B(_2959__bF_buf3), .C(_2961_), .Y(_1661_) );
	OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_24__2_), .Y(_2962_) );
	OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf2), .B(_2959__bF_buf2), .C(_2962_), .Y(_1662_) );
	OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_24__3_), .Y(_2963_) );
	OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf2), .B(_2959__bF_buf1), .C(_2963_), .Y(_1663_) );
	OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_24__4_), .Y(_2964_) );
	OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf2), .B(_2959__bF_buf0), .C(_2964_), .Y(_1664_) );
	OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_24__5_), .Y(_2965_) );
	OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf2), .B(_2959__bF_buf4), .C(_2965_), .Y(_1665_) );
	OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_24__6_), .Y(_2966_) );
	OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf2), .B(_2959__bF_buf3), .C(_2966_), .Y(_1666_) );
	OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_24__7_), .Y(_2967_) );
	OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf2), .B(_2959__bF_buf2), .C(_2967_), .Y(_1667_) );
	OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_24__8_), .Y(_2968_) );
	OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf2), .B(_2959__bF_buf1), .C(_2968_), .Y(_1668_) );
	OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_24__9_), .Y(_2969_) );
	OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf2), .B(_2959__bF_buf0), .C(_2969_), .Y(_1669_) );
	OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_24__10_), .Y(_2970_) );
	OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf2), .B(_2959__bF_buf4), .C(_2970_), .Y(_1670_) );
	OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_24__11_), .Y(_2971_) );
	OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf2), .B(_2959__bF_buf3), .C(_2971_), .Y(_1671_) );
	OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_24__12_), .Y(_2972_) );
	OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf2), .B(_2959__bF_buf2), .C(_2972_), .Y(_1672_) );
	OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_24__13_), .Y(_2973_) );
	OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf2), .B(_2959__bF_buf1), .C(_2973_), .Y(_1673_) );
	OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_24__14_), .Y(_2974_) );
	OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf2), .B(_2959__bF_buf0), .C(_2974_), .Y(_1674_) );
	OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_24__15_), .Y(_2975_) );
	OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf2), .B(_2959__bF_buf4), .C(_2975_), .Y(_1675_) );
	OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_24__16_), .Y(_2976_) );
	OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf2), .B(_2959__bF_buf3), .C(_2976_), .Y(_1676_) );
	OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_24__17_), .Y(_2977_) );
	OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf2), .B(_2959__bF_buf2), .C(_2977_), .Y(_1677_) );
	OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_24__18_), .Y(_2978_) );
	OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf2), .B(_2959__bF_buf1), .C(_2978_), .Y(_1678_) );
	OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_24__19_), .Y(_2979_) );
	OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf2), .B(_2959__bF_buf0), .C(_2979_), .Y(_1679_) );
	OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_24__20_), .Y(_2980_) );
	OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf2), .B(_2959__bF_buf4), .C(_2980_), .Y(_1680_) );
	OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_2553__bF_buf3), .C(csr_gpr_iu_gpr_24__21_), .Y(_2981_) );
	OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf2), .B(_2959__bF_buf3), .C(_2981_), .Y(_1681_) );
	OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_2553__bF_buf2), .C(csr_gpr_iu_gpr_24__22_), .Y(_2982_) );
	OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf2), .B(_2959__bF_buf2), .C(_2982_), .Y(_1682_) );
	OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_2553__bF_buf1), .C(csr_gpr_iu_gpr_24__23_), .Y(_2983_) );
	OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf2), .B(_2959__bF_buf1), .C(_2983_), .Y(_1683_) );
	OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_2553__bF_buf0), .C(csr_gpr_iu_gpr_24__24_), .Y(_2984_) );
	OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf2), .B(_2959__bF_buf0), .C(_2984_), .Y(_1684_) );
	OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_2553__bF_buf10), .C(csr_gpr_iu_gpr_24__25_), .Y(_2985_) );
	OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf2), .B(_2959__bF_buf4), .C(_2985_), .Y(_1685_) );
	OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_2553__bF_buf9), .C(csr_gpr_iu_gpr_24__26_), .Y(_2986_) );
	OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf2), .B(_2959__bF_buf3), .C(_2986_), .Y(_1686_) );
	OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_2553__bF_buf8), .C(csr_gpr_iu_gpr_24__27_), .Y(_2987_) );
	OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf2), .B(_2959__bF_buf2), .C(_2987_), .Y(_1687_) );
	OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_2553__bF_buf7), .C(csr_gpr_iu_gpr_24__28_), .Y(_2988_) );
	OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf2), .B(_2959__bF_buf1), .C(_2988_), .Y(_1688_) );
	OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_2553__bF_buf6), .C(csr_gpr_iu_gpr_24__29_), .Y(_2989_) );
	OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf2), .B(_2959__bF_buf0), .C(_2989_), .Y(_1689_) );
	OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_2553__bF_buf5), .C(csr_gpr_iu_gpr_24__30_), .Y(_2990_) );
	OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_2959__bF_buf4), .C(_2990_), .Y(_1690_) );
	OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_2553__bF_buf4), .C(csr_gpr_iu_gpr_24__31_), .Y(_2991_) );
	OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf2), .B(_2959__bF_buf3), .C(_2991_), .Y(_1691_) );
	INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__0_), .Y(_2992_) );
	NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2479_), .C(_2551_), .Y(_2993_) );
	NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2590__bF_buf12), .Y(_2994_) );
	INVX8 INVX8_46 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .Y(_2995_) );
	NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2995__bF_buf8), .C(_2588__bF_buf5), .Y(_2996_) );
	OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_2994__bF_buf4), .C(_2996_), .Y(_1692_) );
	INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__1_), .Y(_2997_) );
	NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2995__bF_buf7), .C(_2588__bF_buf4), .Y(_2998_) );
	OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_2994__bF_buf3), .C(_2998_), .Y(_1693_) );
	INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__2_), .Y(_2999_) );
	NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2995__bF_buf6), .C(_2588__bF_buf3), .Y(_3000_) );
	OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_2994__bF_buf2), .C(_3000_), .Y(_1694_) );
	INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__3_), .Y(_3001_) );
	NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2995__bF_buf5), .C(_2588__bF_buf2), .Y(_3002_) );
	OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(_2994__bF_buf1), .C(_3002_), .Y(_1695_) );
	INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__4_), .Y(_3003_) );
	NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2995__bF_buf4), .C(_2588__bF_buf1), .Y(_3004_) );
	OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_2994__bF_buf0), .C(_3004_), .Y(_1696_) );
	INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__5_), .Y(_3005_) );
	NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2995__bF_buf3), .C(_2588__bF_buf0), .Y(_3006_) );
	OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_2994__bF_buf4), .C(_3006_), .Y(_1697_) );
	INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__6_), .Y(_3007_) );
	NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2995__bF_buf2), .C(_2588__bF_buf7), .Y(_3008_) );
	OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(_2994__bF_buf3), .C(_3008_), .Y(_1698_) );
	INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__7_), .Y(_3009_) );
	NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2995__bF_buf1), .C(_2588__bF_buf6), .Y(_3010_) );
	OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_2994__bF_buf2), .C(_3010_), .Y(_1699_) );
	INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__8_), .Y(_3011_) );
	NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2995__bF_buf0), .C(_2588__bF_buf5), .Y(_3012_) );
	OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_3011_), .B(_2994__bF_buf1), .C(_3012_), .Y(_1700_) );
	INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__9_), .Y(_3013_) );
	NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2995__bF_buf8), .C(_2588__bF_buf4), .Y(_3014_) );
	OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_2994__bF_buf0), .C(_3014_), .Y(_1701_) );
	INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__10_), .Y(_3015_) );
	NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2995__bF_buf7), .C(_2588__bF_buf3), .Y(_3016_) );
	OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_3015_), .B(_2994__bF_buf4), .C(_3016_), .Y(_1702_) );
	INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__11_), .Y(_3017_) );
	NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2995__bF_buf6), .C(_2588__bF_buf2), .Y(_3018_) );
	OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .B(_2994__bF_buf3), .C(_3018_), .Y(_1703_) );
	INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__12_), .Y(_3019_) );
	NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2995__bF_buf5), .C(_2588__bF_buf1), .Y(_3020_) );
	OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_2994__bF_buf2), .C(_3020_), .Y(_1704_) );
	INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__13_), .Y(_3021_) );
	NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2995__bF_buf4), .C(_2588__bF_buf0), .Y(_3022_) );
	OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_2994__bF_buf1), .C(_3022_), .Y(_1705_) );
	INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__14_), .Y(_3023_) );
	NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2995__bF_buf3), .C(_2588__bF_buf7), .Y(_3024_) );
	OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_2994__bF_buf0), .C(_3024_), .Y(_1706_) );
	INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__15_), .Y(_3025_) );
	NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2995__bF_buf2), .C(_2588__bF_buf6), .Y(_3026_) );
	OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_2994__bF_buf4), .C(_3026_), .Y(_1707_) );
	INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__16_), .Y(_3027_) );
	NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2995__bF_buf1), .C(_2588__bF_buf5), .Y(_3028_) );
	OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_2994__bF_buf3), .C(_3028_), .Y(_1708_) );
	INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__17_), .Y(_3029_) );
	NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2995__bF_buf0), .C(_2588__bF_buf4), .Y(_3030_) );
	OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .B(_2994__bF_buf2), .C(_3030_), .Y(_1709_) );
	INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__18_), .Y(_3031_) );
	NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2995__bF_buf8), .C(_2588__bF_buf3), .Y(_3032_) );
	OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_2994__bF_buf1), .C(_3032_), .Y(_1710_) );
	INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__19_), .Y(_3033_) );
	NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2995__bF_buf7), .C(_2588__bF_buf2), .Y(_3034_) );
	OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .B(_2994__bF_buf0), .C(_3034_), .Y(_1711_) );
	INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__20_), .Y(_3035_) );
	NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2995__bF_buf6), .C(_2588__bF_buf1), .Y(_3036_) );
	OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_2994__bF_buf4), .C(_3036_), .Y(_1712_) );
	INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__21_), .Y(_3037_) );
	NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2995__bF_buf5), .C(_2588__bF_buf0), .Y(_3038_) );
	OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_2994__bF_buf3), .C(_3038_), .Y(_1713_) );
	INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__22_), .Y(_3039_) );
	NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2995__bF_buf4), .C(_2588__bF_buf7), .Y(_3040_) );
	OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .B(_2994__bF_buf2), .C(_3040_), .Y(_1714_) );
	INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__23_), .Y(_3041_) );
	NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2995__bF_buf3), .C(_2588__bF_buf6), .Y(_3042_) );
	OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_2994__bF_buf1), .C(_3042_), .Y(_1715_) );
	INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__24_), .Y(_3043_) );
	NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2995__bF_buf2), .C(_2588__bF_buf5), .Y(_3044_) );
	OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_2994__bF_buf0), .C(_3044_), .Y(_1716_) );
	INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__25_), .Y(_3045_) );
	NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2995__bF_buf1), .C(_2588__bF_buf4), .Y(_3046_) );
	OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_3045_), .B(_2994__bF_buf4), .C(_3046_), .Y(_1717_) );
	INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__26_), .Y(_3047_) );
	NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2995__bF_buf0), .C(_2588__bF_buf3), .Y(_3048_) );
	OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_2994__bF_buf3), .C(_3048_), .Y(_1718_) );
	INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__27_), .Y(_3049_) );
	NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2995__bF_buf8), .C(_2588__bF_buf2), .Y(_3050_) );
	OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_2994__bF_buf2), .C(_3050_), .Y(_1719_) );
	INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__28_), .Y(_3051_) );
	NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2995__bF_buf7), .C(_2588__bF_buf1), .Y(_3052_) );
	OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_2994__bF_buf1), .C(_3052_), .Y(_1720_) );
	INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__29_), .Y(_3053_) );
	NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2995__bF_buf6), .C(_2588__bF_buf0), .Y(_3054_) );
	OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_2994__bF_buf0), .C(_3054_), .Y(_1721_) );
	INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__30_), .Y(_3055_) );
	NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2995__bF_buf5), .C(_2588__bF_buf7), .Y(_3056_) );
	OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_2994__bF_buf4), .C(_3056_), .Y(_1722_) );
	INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_18__31_), .Y(_3057_) );
	NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2995__bF_buf4), .C(_2588__bF_buf6), .Y(_3058_) );
	OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .B(_2994__bF_buf3), .C(_3058_), .Y(_1723_) );
	NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2995__bF_buf3), .B(_2623_), .Y(_3059_) );
	OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf10), .C(csr_gpr_iu_gpr_19__0_), .Y(_3060_) );
	OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf1), .B(_3059__bF_buf4), .C(_3060_), .Y(_1724_) );
	OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf9), .C(csr_gpr_iu_gpr_19__1_), .Y(_3061_) );
	OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf1), .B(_3059__bF_buf3), .C(_3061_), .Y(_1725_) );
	OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2625__bF_buf8), .C(csr_gpr_iu_gpr_19__2_), .Y(_3062_) );
	OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf1), .B(_3059__bF_buf2), .C(_3062_), .Y(_1726_) );
	OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2625__bF_buf7), .C(csr_gpr_iu_gpr_19__3_), .Y(_3063_) );
	OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf1), .B(_3059__bF_buf1), .C(_3063_), .Y(_1727_) );
	OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2625__bF_buf6), .C(csr_gpr_iu_gpr_19__4_), .Y(_3064_) );
	OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf1), .B(_3059__bF_buf0), .C(_3064_), .Y(_1728_) );
	OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .B(_2625__bF_buf5), .C(csr_gpr_iu_gpr_19__5_), .Y(_3065_) );
	OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf1), .B(_3059__bF_buf4), .C(_3065_), .Y(_1729_) );
	OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf4), .C(csr_gpr_iu_gpr_19__6_), .Y(_3066_) );
	OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf1), .B(_3059__bF_buf3), .C(_3066_), .Y(_1730_) );
	OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf3), .C(csr_gpr_iu_gpr_19__7_), .Y(_3067_) );
	OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf1), .B(_3059__bF_buf2), .C(_3067_), .Y(_1731_) );
	OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2625__bF_buf2), .C(csr_gpr_iu_gpr_19__8_), .Y(_3068_) );
	OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf1), .B(_3059__bF_buf1), .C(_3068_), .Y(_1732_) );
	OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2625__bF_buf1), .C(csr_gpr_iu_gpr_19__9_), .Y(_3069_) );
	OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf1), .B(_3059__bF_buf0), .C(_3069_), .Y(_1733_) );
	OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2625__bF_buf0), .C(csr_gpr_iu_gpr_19__10_), .Y(_3070_) );
	OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf1), .B(_3059__bF_buf4), .C(_3070_), .Y(_1734_) );
	OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .B(_2625__bF_buf14), .C(csr_gpr_iu_gpr_19__11_), .Y(_3071_) );
	OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf1), .B(_3059__bF_buf3), .C(_3071_), .Y(_1735_) );
	OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf13), .C(csr_gpr_iu_gpr_19__12_), .Y(_3072_) );
	OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf1), .B(_3059__bF_buf2), .C(_3072_), .Y(_1736_) );
	OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf12), .C(csr_gpr_iu_gpr_19__13_), .Y(_3073_) );
	OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf1), .B(_3059__bF_buf1), .C(_3073_), .Y(_1737_) );
	OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2625__bF_buf11), .C(csr_gpr_iu_gpr_19__14_), .Y(_3074_) );
	OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf1), .B(_3059__bF_buf0), .C(_3074_), .Y(_1738_) );
	OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2625__bF_buf10), .C(csr_gpr_iu_gpr_19__15_), .Y(_3075_) );
	OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf1), .B(_3059__bF_buf4), .C(_3075_), .Y(_1739_) );
	OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2625__bF_buf9), .C(csr_gpr_iu_gpr_19__16_), .Y(_3076_) );
	OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf1), .B(_3059__bF_buf3), .C(_3076_), .Y(_1740_) );
	OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .B(_2625__bF_buf8), .C(csr_gpr_iu_gpr_19__17_), .Y(_3077_) );
	OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf1), .B(_3059__bF_buf2), .C(_3077_), .Y(_1741_) );
	OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf7), .C(csr_gpr_iu_gpr_19__18_), .Y(_3078_) );
	OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf1), .B(_3059__bF_buf1), .C(_3078_), .Y(_1742_) );
	OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf6), .C(csr_gpr_iu_gpr_19__19_), .Y(_3079_) );
	OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf1), .B(_3059__bF_buf0), .C(_3079_), .Y(_1743_) );
	OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2625__bF_buf5), .C(csr_gpr_iu_gpr_19__20_), .Y(_3080_) );
	OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf1), .B(_3059__bF_buf4), .C(_3080_), .Y(_1744_) );
	OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2625__bF_buf4), .C(csr_gpr_iu_gpr_19__21_), .Y(_3081_) );
	OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf1), .B(_3059__bF_buf3), .C(_3081_), .Y(_1745_) );
	OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2625__bF_buf3), .C(csr_gpr_iu_gpr_19__22_), .Y(_3082_) );
	OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf1), .B(_3059__bF_buf2), .C(_3082_), .Y(_1746_) );
	OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .B(_2625__bF_buf2), .C(csr_gpr_iu_gpr_19__23_), .Y(_3083_) );
	OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf1), .B(_3059__bF_buf1), .C(_3083_), .Y(_1747_) );
	OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf1), .C(csr_gpr_iu_gpr_19__24_), .Y(_3084_) );
	OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf1), .B(_3059__bF_buf0), .C(_3084_), .Y(_1748_) );
	OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf0), .C(csr_gpr_iu_gpr_19__25_), .Y(_3085_) );
	OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf1), .B(_3059__bF_buf4), .C(_3085_), .Y(_1749_) );
	OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2625__bF_buf14), .C(csr_gpr_iu_gpr_19__26_), .Y(_3086_) );
	OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf1), .B(_3059__bF_buf3), .C(_3086_), .Y(_1750_) );
	OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2625__bF_buf13), .C(csr_gpr_iu_gpr_19__27_), .Y(_3087_) );
	OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf1), .B(_3059__bF_buf2), .C(_3087_), .Y(_1751_) );
	OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf5), .B(_2625__bF_buf12), .C(csr_gpr_iu_gpr_19__28_), .Y(_3088_) );
	OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf1), .B(_3059__bF_buf1), .C(_3088_), .Y(_1752_) );
	OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf4), .B(_2625__bF_buf11), .C(csr_gpr_iu_gpr_19__29_), .Y(_3089_) );
	OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf1), .B(_3059__bF_buf0), .C(_3089_), .Y(_1753_) );
	OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf3), .B(_2625__bF_buf10), .C(csr_gpr_iu_gpr_19__30_), .Y(_3090_) );
	OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_3059__bF_buf4), .C(_3090_), .Y(_1754_) );
	OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf2), .B(_2625__bF_buf9), .C(csr_gpr_iu_gpr_19__31_), .Y(_3091_) );
	OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf1), .B(_3059__bF_buf3), .C(_3091_), .Y(_1755_) );
	INVX8 INVX8_47 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_19_), .Y(_3092_) );
	INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_17_), .Y(_3093_) );
	INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .Y(_3094_) );
	NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf5), .B(biu_ins_16_), .Y(_3095_) );
	NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_3094_), .C(_3095__bF_buf11), .Y(_3096_) );
	INVX8 INVX8_48 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .Y(_3097_) );
	NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .Y(_3098_) );
	NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_3095__bF_buf10), .Y(_3099_) );
	OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .B(_3099_), .C(biu_ins_19_), .Y(_3100_) );
	NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf3), .B(_3098_), .Y(_3101_) );
	OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_3099_), .B(_3094_), .Y(_3102_) );
	INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf4), .Y(_3103_) );
	INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_16_), .Y(_3104_) );
	NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(_3104_), .Y(_3105_) );
	OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_17_), .B(_3105__bF_buf7), .C(_3094_), .Y(_3106_) );
	NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .B(_3102_), .Y(_3107_) );
	OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf3), .B(biu_ins_16_), .C(biu_ins_17_), .Y(_3108_) );
	NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .B(_3099_), .Y(_3109_) );
	NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf2), .B(biu_ins_16_), .Y(_3110_) );
	NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_16_), .B(_3103_), .Y(_3111_) );
	OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_3110__bF_buf13), .C(_2796_), .D(_3111__bF_buf15), .Y(_3112_) );
	NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf1), .B(_3104_), .Y(_3113_) );
	NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__0_), .B(_3095__bF_buf9), .Y(_3114_) );
	OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_2729_), .B(_3113__bF_buf15), .C(_3114_), .Y(_3115_) );
	OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_3112_), .B(_3115_), .C(_3109__bF_buf10), .Y(_3116_) );
	AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_3099_), .B(_3108_), .Y(_3117_) );
	INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__0_), .Y(_3118_) );
	OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_3110__bF_buf12), .C(_3118_), .D(_3111__bF_buf14), .Y(_3119_) );
	INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__0_), .Y(_3120_) );
	NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__0_), .B(_3095__bF_buf8), .Y(_3121_) );
	OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_3113__bF_buf14), .C(_3121_), .Y(_3122_) );
	OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_3119_), .B(_3122_), .C(_3117__bF_buf9), .Y(_3123_) );
	NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_3116_), .B(_3123_), .C(_3107__bF_buf5), .Y(_3124_) );
	OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_17_), .B(_3105__bF_buf6), .C(biu_ins_18_), .Y(_3125_) );
	NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3125_), .Y(_3126_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf0), .B(biu_ins_16_), .Y(_3127_) );
	NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__0_), .B(_3113__bF_buf13), .C(_3111__bF_buf13), .Y(_3128_) );
	MUX2X1 MUX2X1_59 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__0_), .B(csr_gpr_iu_gpr_29__0_), .S(biu_ins_15_bF_buf6), .Y(_3129_) );
	OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .B(_3127__bF_buf5), .C(_3128_), .Y(_3130_) );
	NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf9), .B(_3130_), .Y(_3131_) );
	INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__0_), .Y(_3132_) );
	NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__0_), .B(_3095__bF_buf7), .Y(_3133_) );
	OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_3132_), .B(_3113__bF_buf12), .C(_3133_), .Y(_3134_) );
	INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__0_), .Y(_3135_) );
	INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__0_), .Y(_3136_) );
	OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3110__bF_buf11), .C(_3135_), .D(_3111__bF_buf12), .Y(_3137_) );
	OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_3137_), .B(_3134_), .C(_3117__bF_buf8), .Y(_3138_) );
	NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf7), .B(_3138_), .C(_3131_), .Y(_3139_) );
	NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3124_), .C(_3139_), .Y(_3140_) );
	INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__0_), .Y(_3141_) );
	INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__0_), .Y(_3142_) );
	OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3142_), .B(_3110__bF_buf10), .C(_3141_), .D(_3113__bF_buf11), .Y(_3143_) );
	INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__0_), .Y(_3144_) );
	NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__0_), .B(_3095__bF_buf6), .Y(_3145_) );
	OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_3111__bF_buf11), .C(_3145_), .Y(_3146_) );
	OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_3146_), .C(_3109__bF_buf8), .Y(_3147_) );
	INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__0_), .Y(_3148_) );
	INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__0_), .Y(_3149_) );
	OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_3110__bF_buf9), .C(_3148_), .D(_3111__bF_buf10), .Y(_3150_) );
	INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__0_), .Y(_3151_) );
	NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__0_), .B(_3095__bF_buf5), .Y(_3152_) );
	OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_3151_), .B(_3113__bF_buf10), .C(_3152_), .Y(_3153_) );
	OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .B(_3153_), .C(_3117__bF_buf7), .Y(_3154_) );
	AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3125_), .C(_3147_), .D(_3154_), .Y(_3155_) );
	INVX8 INVX8_49 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .Y(_3156_) );
	INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__0_), .Y(_3157_) );
	NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__0_), .B(_3095__bF_buf4), .Y(_3158_) );
	OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .B(_3113__bF_buf9), .C(_3158_), .Y(_3159_) );
	INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__0_), .Y(_3160_) );
	INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__0_), .Y(_3161_) );
	OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3110__bF_buf8), .C(_3160_), .D(_3111__bF_buf9), .Y(_3162_) );
	OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .B(_3159_), .C(_3109__bF_buf7), .Y(_3163_) );
	INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__0_), .Y(_3164_) );
	NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__0_), .B(_3095__bF_buf3), .Y(_3165_) );
	OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_3164_), .B(_3113__bF_buf8), .C(_3165_), .Y(_3166_) );
	INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__0_), .Y(_3167_) );
	INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__0_), .Y(_3168_) );
	OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3168_), .B(_3110__bF_buf7), .C(_3167_), .D(_3111__bF_buf8), .Y(_3169_) );
	OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_3166_), .C(_3117__bF_buf6), .Y(_3170_) );
	AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3163_), .B(_3170_), .C(_3126__bF_buf6), .Y(_3171_) );
	OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_3171_), .C(_3156__bF_buf4), .Y(_3172_) );
	AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3140_), .D(_3172_), .Y(csr_gpr_iu_rs1_0_) );
	NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__1_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_3173_) );
	MUX2X1 MUX2X1_60 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__1_), .B(csr_gpr_iu_gpr_29__1_), .S(biu_ins_15_bF_buf5), .Y(_3174_) );
	OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .B(_3127__bF_buf4), .C(_3173_), .Y(_3175_) );
	NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf6), .B(_3175_), .Y(_3176_) );
	INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__1_), .Y(_3177_) );
	NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__1_), .B(_3095__bF_buf2), .Y(_3178_) );
	OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3113__bF_buf6), .C(_3178_), .Y(_3179_) );
	INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__1_), .Y(_3180_) );
	INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__1_), .Y(_3181_) );
	OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3181_), .B(_3110__bF_buf6), .C(_3180_), .D(_3111__bF_buf6), .Y(_3182_) );
	OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_3182_), .B(_3179_), .C(_3117__bF_buf5), .Y(_3183_) );
	NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf5), .B(_3183_), .C(_3176_), .Y(_3184_) );
	OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_3110__bF_buf5), .C(_2799_), .D(_3111__bF_buf5), .Y(_3185_) );
	NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__1_), .B(_3095__bF_buf1), .Y(_3186_) );
	OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_3113__bF_buf5), .C(_3186_), .Y(_3187_) );
	OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .B(_3187_), .C(_3109__bF_buf5), .Y(_3188_) );
	INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__1_), .Y(_3189_) );
	OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_3110__bF_buf4), .C(_3189_), .D(_3111__bF_buf4), .Y(_3190_) );
	INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__1_), .Y(_3191_) );
	NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__1_), .B(_3095__bF_buf0), .Y(_3192_) );
	OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .B(_3113__bF_buf4), .C(_3192_), .Y(_3193_) );
	OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_3190_), .B(_3193_), .C(_3117__bF_buf4), .Y(_3194_) );
	NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_3188_), .B(_3194_), .C(_3107__bF_buf4), .Y(_3195_) );
	NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3195_), .C(_3184_), .Y(_3196_) );
	INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__1_), .Y(_3197_) );
	INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__1_), .Y(_3198_) );
	OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_3110__bF_buf3), .C(_3197_), .D(_3111__bF_buf3), .Y(_3199_) );
	INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__1_), .Y(_3200_) );
	NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__1_), .B(_3095__bF_buf11), .Y(_3201_) );
	OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(_3113__bF_buf3), .C(_3201_), .Y(_3202_) );
	OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3202_), .C(_3109__bF_buf4), .Y(_3203_) );
	INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__1_), .Y(_3204_) );
	INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__1_), .Y(_3205_) );
	OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3205_), .B(_3110__bF_buf2), .C(_3204_), .D(_3113__bF_buf2), .Y(_3206_) );
	INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__1_), .Y(_3207_) );
	NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__1_), .B(_3095__bF_buf10), .Y(_3208_) );
	OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .B(_3111__bF_buf2), .C(_3208_), .Y(_3209_) );
	OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_3206_), .B(_3209_), .C(_3117__bF_buf3), .Y(_3210_) );
	AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3203_), .D(_3210_), .Y(_3211_) );
	INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__1_), .Y(_3212_) );
	INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__1_), .Y(_3213_) );
	OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3110__bF_buf1), .C(_3212_), .D(_3111__bF_buf1), .Y(_3214_) );
	INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__1_), .Y(_3215_) );
	NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__1_), .B(_3095__bF_buf9), .Y(_3216_) );
	OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3113__bF_buf1), .C(_3216_), .Y(_3217_) );
	OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_3217_), .C(_3109__bF_buf3), .Y(_3218_) );
	INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__1_), .Y(_3219_) );
	INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__1_), .Y(_3220_) );
	OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_3220_), .B(_3110__bF_buf0), .C(_3219_), .D(_3111__bF_buf0), .Y(_3221_) );
	INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__1_), .Y(_3222_) );
	NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__1_), .B(_3095__bF_buf8), .Y(_3223_) );
	OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_3113__bF_buf0), .C(_3223_), .Y(_3224_) );
	OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_3221_), .B(_3224_), .C(_3117__bF_buf2), .Y(_3225_) );
	AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3218_), .B(_3225_), .C(_3107__bF_buf3), .Y(_3226_) );
	OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_3211_), .B(_3226_), .C(_3156__bF_buf3), .Y(_3227_) );
	AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3196_), .D(_3227_), .Y(csr_gpr_iu_rs1_1_) );
	INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__2_), .Y(_3228_) );
	INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__2_), .Y(_3229_) );
	OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_3229_), .B(_3110__bF_buf13), .C(_3228_), .D(_3105__bF_buf5), .Y(_3230_) );
	INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__2_), .Y(_3231_) );
	INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__2_), .Y(_3232_) );
	OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3111__bF_buf15), .C(_3232_), .D(_3113__bF_buf15), .Y(_3233_) );
	OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_3233_), .C(_3109__bF_buf2), .Y(_3234_) );
	INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__2_), .Y(_3235_) );
	INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__2_), .Y(_3236_) );
	OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_3110__bF_buf12), .C(_3235_), .D(_3105__bF_buf4), .Y(_3237_) );
	INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__2_), .Y(_3238_) );
	INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__2_), .Y(_3239_) );
	OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_3111__bF_buf14), .C(_3239_), .D(_3113__bF_buf14), .Y(_3240_) );
	OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_3237_), .B(_3240_), .C(_3117__bF_buf1), .Y(_3241_) );
	AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_3241_), .B(_3234_), .C(_3107__bF_buf2), .Y(_3242_) );
	INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__2_), .Y(_3243_) );
	INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__2_), .Y(_3244_) );
	OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3111__bF_buf13), .C(_3244_), .D(_3113__bF_buf13), .Y(_3245_) );
	INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__2_), .Y(_3246_) );
	NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__2_), .B(_3095__bF_buf7), .Y(_3247_) );
	OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_3110__bF_buf11), .C(_3247_), .Y(_3248_) );
	OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_3245_), .B(_3248_), .C(_3109__bF_buf1), .Y(_3249_) );
	INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__2_), .Y(_3250_) );
	INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__2_), .Y(_3251_) );
	OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_3111__bF_buf12), .C(_3251_), .D(_3113__bF_buf12), .Y(_3252_) );
	INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__2_), .Y(_3253_) );
	NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__2_), .B(_3095__bF_buf6), .Y(_3254_) );
	OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3110__bF_buf10), .C(_3254_), .Y(_3255_) );
	OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .B(_3255_), .C(_3117__bF_buf0), .Y(_3256_) );
	AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_3256_), .C(_3126__bF_buf4), .Y(_3257_) );
	OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .B(_3257_), .C(_3156__bF_buf2), .Y(_3258_) );
	INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__2_), .Y(_3259_) );
	INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__2_), .Y(_3260_) );
	OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_3111__bF_buf11), .C(_3260_), .D(_3113__bF_buf11), .Y(_3261_) );
	INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__2_), .Y(_3262_) );
	NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__2_), .B(biu_ins_15_bF_buf4), .Y(_3263_) );
	OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf3), .B(_3262_), .C(_3263_), .Y(_3264_) );
	AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf3), .B(_3264_), .C(_3261_), .Y(_3265_) );
	INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__2_), .Y(_3266_) );
	INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__2_), .Y(_3267_) );
	OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .B(_3111__bF_buf10), .C(_3267_), .D(_3113__bF_buf10), .Y(_3268_) );
	AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__2_), .B(_3127__bF_buf2), .C(_3268_), .Y(_3269_) );
	MUX2X1 MUX2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3265_), .S(_3109__bF_buf0), .Y(_3270_) );
	NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__2_), .B(_3095__bF_buf5), .Y(_3271_) );
	OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_2801_), .B(_3111__bF_buf9), .C(_3271_), .Y(_3272_) );
	OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_3110__bF_buf9), .C(_2736_), .D(_3113__bF_buf9), .Y(_3273_) );
	OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_3273_), .B(_3272_), .C(_3109__bF_buf10), .Y(_3274_) );
	INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__2_), .Y(_3275_) );
	INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__2_), .Y(_3276_) );
	OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_3111__bF_buf8), .C(_3276_), .D(_3113__bF_buf8), .Y(_3277_) );
	INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__2_), .Y(_3278_) );
	OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_3110__bF_buf8), .C(_3278_), .D(_3105__bF_buf3), .Y(_3279_) );
	OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_3279_), .B(_3277_), .C(_3117__bF_buf9), .Y(_3280_) );
	AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_3280_), .C(_3126__bF_buf3), .Y(_3281_) );
	AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3126__bF_buf2), .C(_3281_), .Y(_3282_) );
	OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf2), .B(_3282_), .C(_3258_), .Y(csr_gpr_iu_rs1_2_) );
	INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__3_), .Y(_3283_) );
	INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__3_), .Y(_3284_) );
	OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_3110__bF_buf7), .C(_3283_), .D(_3105__bF_buf2), .Y(_3285_) );
	INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__3_), .Y(_3286_) );
	INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__3_), .Y(_3287_) );
	OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3111__bF_buf7), .C(_3287_), .D(_3113__bF_buf7), .Y(_3288_) );
	OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_3285_), .B(_3288_), .C(_3109__bF_buf9), .Y(_3289_) );
	INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__3_), .Y(_3290_) );
	INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__3_), .Y(_3291_) );
	OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_3291_), .B(_3110__bF_buf6), .C(_3290_), .D(_3105__bF_buf1), .Y(_3292_) );
	INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__3_), .Y(_3293_) );
	INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__3_), .Y(_3294_) );
	OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_3111__bF_buf6), .C(_3294_), .D(_3113__bF_buf6), .Y(_3295_) );
	OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3295_), .C(_3117__bF_buf8), .Y(_3296_) );
	AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_3289_), .C(_3107__bF_buf1), .Y(_3297_) );
	INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__3_), .Y(_3298_) );
	INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__3_), .Y(_3299_) );
	OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_3110__bF_buf5), .C(_3298_), .D(_3113__bF_buf5), .Y(_3300_) );
	INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__3_), .Y(_3301_) );
	INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__3_), .Y(_3302_) );
	OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_3301_), .B(_3111__bF_buf5), .C(_3302_), .D(_3105__bF_buf0), .Y(_3303_) );
	OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_3300_), .B(_3303_), .C(_3109__bF_buf8), .Y(_3304_) );
	INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__3_), .Y(_3305_) );
	INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__3_), .Y(_3306_) );
	OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_3110__bF_buf4), .C(_3305_), .D(_3113__bF_buf4), .Y(_3307_) );
	INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__3_), .Y(_3308_) );
	INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__3_), .Y(_3309_) );
	OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3111__bF_buf4), .C(_3309_), .D(_3105__bF_buf7), .Y(_3310_) );
	OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_3310_), .C(_3117__bF_buf7), .Y(_3311_) );
	AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_3304_), .C(_3126__bF_buf1), .Y(_3312_) );
	OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_3297_), .B(_3312_), .C(_3156__bF_buf1), .Y(_3313_) );
	INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__3_), .Y(_3314_) );
	INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__3_), .Y(_3315_) );
	OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_3111__bF_buf3), .C(_3315_), .D(_3113__bF_buf3), .Y(_3316_) );
	INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__3_), .Y(_3317_) );
	NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__3_), .B(biu_ins_15_bF_buf2), .Y(_3318_) );
	OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf1), .B(_3317_), .C(_3318_), .Y(_3319_) );
	AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf1), .B(_3319_), .C(_3316_), .Y(_3320_) );
	INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__3_), .Y(_3321_) );
	INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__3_), .Y(_3322_) );
	OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(_3111__bF_buf2), .C(_3322_), .D(_3113__bF_buf2), .Y(_3323_) );
	AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__3_), .B(_3127__bF_buf0), .C(_3323_), .Y(_3324_) );
	MUX2X1 MUX2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_3320_), .S(_3109__bF_buf7), .Y(_3325_) );
	NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__3_), .B(_3095__bF_buf4), .Y(_3326_) );
	OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_3111__bF_buf1), .C(_3326_), .Y(_3327_) );
	OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(_3110__bF_buf3), .C(_2738_), .D(_3113__bF_buf1), .Y(_3328_) );
	OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3327_), .C(_3109__bF_buf6), .Y(_3329_) );
	INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__3_), .Y(_3330_) );
	INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__3_), .Y(_3331_) );
	OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_3111__bF_buf0), .C(_3331_), .D(_3113__bF_buf0), .Y(_3332_) );
	INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__3_), .Y(_3333_) );
	OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(_3110__bF_buf2), .C(_3333_), .D(_3105__bF_buf6), .Y(_3334_) );
	OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_3334_), .B(_3332_), .C(_3117__bF_buf6), .Y(_3335_) );
	AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3335_), .C(_3126__bF_buf0), .Y(_3336_) );
	AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_3126__bF_buf7), .C(_3336_), .Y(_3337_) );
	OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf1), .B(_3337_), .C(_3313_), .Y(csr_gpr_iu_rs1_3_) );
	NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__4_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_3338_) );
	MUX2X1 MUX2X1_63 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__4_), .B(csr_gpr_iu_gpr_29__4_), .S(biu_ins_15_bF_buf0), .Y(_3339_) );
	OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_3127__bF_buf5), .C(_3338_), .Y(_3340_) );
	NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf5), .B(_3340_), .Y(_3341_) );
	INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__4_), .Y(_3342_) );
	NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__4_), .B(_3095__bF_buf3), .Y(_3343_) );
	OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .B(_3113__bF_buf14), .C(_3343_), .Y(_3344_) );
	INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__4_), .Y(_3345_) );
	INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__4_), .Y(_3346_) );
	OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3110__bF_buf1), .C(_3345_), .D(_3111__bF_buf14), .Y(_3347_) );
	OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_3347_), .B(_3344_), .C(_3117__bF_buf5), .Y(_3348_) );
	NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf6), .B(_3348_), .C(_3341_), .Y(_3349_) );
	NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__4_), .B(_3095__bF_buf2), .Y(_3350_) );
	OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_3111__bF_buf13), .C(_3350_), .Y(_3351_) );
	OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_3110__bF_buf0), .C(_2740_), .D(_3113__bF_buf13), .Y(_3352_) );
	OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .B(_3351_), .C(_3109__bF_buf4), .Y(_3353_) );
	INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__4_), .Y(_3354_) );
	NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__4_), .B(_3095__bF_buf1), .Y(_3355_) );
	OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(_3111__bF_buf12), .C(_3355_), .Y(_3356_) );
	INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__4_), .Y(_3357_) );
	OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_3110__bF_buf13), .C(_3357_), .D(_3113__bF_buf12), .Y(_3358_) );
	OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_3358_), .B(_3356_), .C(_3117__bF_buf4), .Y(_3359_) );
	NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .B(_3359_), .C(_3107__bF_buf0), .Y(_3360_) );
	NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3360_), .C(_3349_), .Y(_3361_) );
	INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__4_), .Y(_3362_) );
	NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__4_), .B(_3095__bF_buf0), .Y(_3363_) );
	OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3111__bF_buf11), .C(_3363_), .Y(_3364_) );
	INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__4_), .Y(_3365_) );
	INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__4_), .Y(_3366_) );
	OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_3110__bF_buf12), .C(_3365_), .D(_3113__bF_buf11), .Y(_3367_) );
	OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_3364_), .C(_3109__bF_buf3), .Y(_3368_) );
	INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__4_), .Y(_3369_) );
	NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__4_), .B(_3095__bF_buf11), .Y(_3370_) );
	OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_3113__bF_buf10), .C(_3370_), .Y(_3371_) );
	INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__4_), .Y(_3372_) );
	INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__4_), .Y(_3373_) );
	OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3110__bF_buf11), .C(_3372_), .D(_3111__bF_buf10), .Y(_3374_) );
	OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3371_), .C(_3117__bF_buf3), .Y(_3375_) );
	AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3368_), .D(_3375_), .Y(_3376_) );
	INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__4_), .Y(_3377_) );
	NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__4_), .B(_3095__bF_buf10), .Y(_3378_) );
	OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_3377_), .B(_3111__bF_buf9), .C(_3378_), .Y(_3379_) );
	INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__4_), .Y(_3380_) );
	INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__4_), .Y(_3381_) );
	OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3110__bF_buf10), .C(_3380_), .D(_3113__bF_buf9), .Y(_3382_) );
	OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3379_), .C(_3109__bF_buf2), .Y(_3383_) );
	INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__4_), .Y(_3384_) );
	NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__4_), .B(_3095__bF_buf9), .Y(_3385_) );
	OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3111__bF_buf8), .C(_3385_), .Y(_3386_) );
	INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__4_), .Y(_3387_) );
	INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__4_), .Y(_3388_) );
	OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3110__bF_buf9), .C(_3387_), .D(_3113__bF_buf8), .Y(_3389_) );
	OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3386_), .C(_3117__bF_buf2), .Y(_3390_) );
	AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3383_), .B(_3390_), .C(_3107__bF_buf5), .Y(_3391_) );
	OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .B(_3391_), .C(_3156__bF_buf0), .Y(_3392_) );
	AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3361_), .D(_3392_), .Y(csr_gpr_iu_rs1_4_) );
	INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__5_), .Y(_3393_) );
	INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__5_), .Y(_3394_) );
	OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3394_), .B(_3110__bF_buf8), .C(_3393_), .D(_3105__bF_buf5), .Y(_3395_) );
	INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__5_), .Y(_3396_) );
	INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__5_), .Y(_3397_) );
	OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_3111__bF_buf7), .C(_3397_), .D(_3113__bF_buf7), .Y(_3398_) );
	OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .B(_3398_), .C(_3109__bF_buf1), .Y(_3399_) );
	INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__5_), .Y(_3400_) );
	INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__5_), .Y(_3401_) );
	OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3401_), .B(_3110__bF_buf7), .C(_3400_), .D(_3105__bF_buf4), .Y(_3402_) );
	INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__5_), .Y(_3403_) );
	INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__5_), .Y(_3404_) );
	OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_3111__bF_buf6), .C(_3404_), .D(_3113__bF_buf6), .Y(_3405_) );
	OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3405_), .C(_3117__bF_buf1), .Y(_3406_) );
	AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3399_), .C(_3107__bF_buf4), .Y(_3407_) );
	INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__5_), .Y(_3408_) );
	NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__5_), .B(_3095__bF_buf8), .Y(_3409_) );
	OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3113__bF_buf5), .C(_3409_), .Y(_3410_) );
	INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__5_), .Y(_3411_) );
	INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__5_), .Y(_3412_) );
	OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3110__bF_buf6), .C(_3411_), .D(_3111__bF_buf5), .Y(_3413_) );
	OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_3410_), .C(_3109__bF_buf0), .Y(_3414_) );
	INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__5_), .Y(_3415_) );
	NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__5_), .B(_3095__bF_buf7), .Y(_3416_) );
	OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_3415_), .B(_3113__bF_buf4), .C(_3416_), .Y(_3417_) );
	INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__5_), .Y(_3418_) );
	INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__5_), .Y(_3419_) );
	OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3110__bF_buf5), .C(_3418_), .D(_3111__bF_buf4), .Y(_3420_) );
	OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .B(_3417_), .C(_3117__bF_buf0), .Y(_3421_) );
	AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3414_), .B(_3421_), .C(_3126__bF_buf5), .Y(_3422_) );
	OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_3407_), .B(_3422_), .C(_3156__bF_buf4), .Y(_3423_) );
	INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__5_), .Y(_3424_) );
	INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__5_), .Y(_3425_) );
	OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3424_), .B(_3111__bF_buf3), .C(_3425_), .D(_3113__bF_buf3), .Y(_3426_) );
	INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__5_), .Y(_3427_) );
	NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__5_), .B(biu_ins_15_bF_buf6), .Y(_3428_) );
	OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf5), .B(_3427_), .C(_3428_), .Y(_3429_) );
	AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf4), .B(_3429_), .C(_3426_), .Y(_3430_) );
	INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__5_), .Y(_3431_) );
	INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__5_), .Y(_3432_) );
	OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .B(_3111__bF_buf2), .C(_3432_), .D(_3113__bF_buf2), .Y(_3433_) );
	AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__5_), .B(_3127__bF_buf3), .C(_3433_), .Y(_3434_) );
	MUX2X1 MUX2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .B(_3430_), .S(_3109__bF_buf10), .Y(_3435_) );
	OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_3110__bF_buf4), .C(_2807_), .D(_3111__bF_buf1), .Y(_3436_) );
	NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__5_), .B(_3095__bF_buf6), .Y(_3437_) );
	OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_3113__bF_buf1), .C(_3437_), .Y(_3438_) );
	OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_3436_), .B(_3438_), .C(_3109__bF_buf9), .Y(_3439_) );
	INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__5_), .Y(_3440_) );
	INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__5_), .Y(_3441_) );
	OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_3111__bF_buf0), .C(_3441_), .D(_3113__bF_buf0), .Y(_3442_) );
	INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__5_), .Y(_3443_) );
	OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_3110__bF_buf3), .C(_3443_), .D(_3105__bF_buf3), .Y(_3444_) );
	OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_3444_), .B(_3442_), .C(_3117__bF_buf9), .Y(_3445_) );
	AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3445_), .C(_3126__bF_buf4), .Y(_3446_) );
	AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .B(_3126__bF_buf3), .C(_3446_), .Y(_3447_) );
	OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf0), .B(_3447_), .C(_3423_), .Y(csr_gpr_iu_rs1_5_) );
	INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__6_), .Y(_3448_) );
	INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__6_), .Y(_3449_) );
	OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3110__bF_buf2), .C(_3448_), .D(_3105__bF_buf2), .Y(_3450_) );
	INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__6_), .Y(_3451_) );
	INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__6_), .Y(_3452_) );
	OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_3111__bF_buf15), .C(_3452_), .D(_3113__bF_buf15), .Y(_3453_) );
	OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_3450_), .B(_3453_), .C(_3109__bF_buf8), .Y(_3454_) );
	INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__6_), .Y(_3455_) );
	INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__6_), .Y(_3456_) );
	OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3456_), .B(_3110__bF_buf1), .C(_3455_), .D(_3105__bF_buf1), .Y(_3457_) );
	INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__6_), .Y(_3458_) );
	INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__6_), .Y(_3459_) );
	OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3111__bF_buf14), .C(_3459_), .D(_3113__bF_buf14), .Y(_3460_) );
	OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_3460_), .C(_3117__bF_buf8), .Y(_3461_) );
	AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .B(_3454_), .C(_3107__bF_buf3), .Y(_3462_) );
	INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__6_), .Y(_3463_) );
	NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__6_), .B(_3095__bF_buf5), .Y(_3464_) );
	OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_3463_), .B(_3113__bF_buf13), .C(_3464_), .Y(_3465_) );
	INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__6_), .Y(_3466_) );
	INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__6_), .Y(_3467_) );
	OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3110__bF_buf0), .C(_3466_), .D(_3111__bF_buf13), .Y(_3468_) );
	OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_3468_), .B(_3465_), .C(_3109__bF_buf7), .Y(_3469_) );
	INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__6_), .Y(_3470_) );
	NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__6_), .B(_3095__bF_buf4), .Y(_3471_) );
	OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3113__bF_buf12), .C(_3471_), .Y(_3472_) );
	INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__6_), .Y(_3473_) );
	INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__6_), .Y(_3474_) );
	OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(_3110__bF_buf13), .C(_3473_), .D(_3111__bF_buf12), .Y(_3475_) );
	OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_3475_), .B(_3472_), .C(_3117__bF_buf7), .Y(_3476_) );
	AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3476_), .C(_3126__bF_buf2), .Y(_3477_) );
	OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3477_), .C(_3156__bF_buf3), .Y(_3478_) );
	INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__6_), .Y(_3479_) );
	INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__6_), .Y(_3480_) );
	OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_3111__bF_buf11), .C(_3480_), .D(_3113__bF_buf11), .Y(_3481_) );
	INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__6_), .Y(_3482_) );
	NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__6_), .B(biu_ins_15_bF_buf4), .Y(_3483_) );
	OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf3), .B(_3482_), .C(_3483_), .Y(_3484_) );
	AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf2), .B(_3484_), .C(_3481_), .Y(_3485_) );
	INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__6_), .Y(_3486_) );
	INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__6_), .Y(_3487_) );
	OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_3111__bF_buf10), .C(_3487_), .D(_3113__bF_buf10), .Y(_3488_) );
	AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__6_), .B(_3127__bF_buf1), .C(_3488_), .Y(_3489_) );
	MUX2X1 MUX2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_3485_), .S(_3109__bF_buf6), .Y(_3490_) );
	NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__6_), .B(_3095__bF_buf3), .Y(_3491_) );
	OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_2809_), .B(_3111__bF_buf9), .C(_3491_), .Y(_3492_) );
	OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .B(_3110__bF_buf12), .C(_2744_), .D(_3113__bF_buf9), .Y(_3493_) );
	OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_3493_), .B(_3492_), .C(_3109__bF_buf5), .Y(_3494_) );
	INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__6_), .Y(_3495_) );
	INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__6_), .Y(_3496_) );
	OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_3111__bF_buf8), .C(_3496_), .D(_3113__bF_buf8), .Y(_3497_) );
	INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__6_), .Y(_3498_) );
	OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(_3110__bF_buf11), .C(_3498_), .D(_3105__bF_buf0), .Y(_3499_) );
	OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_3497_), .C(_3117__bF_buf6), .Y(_3500_) );
	AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .B(_3500_), .C(_3126__bF_buf1), .Y(_3501_) );
	AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(_3126__bF_buf0), .C(_3501_), .Y(_3502_) );
	OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf3), .B(_3502_), .C(_3478_), .Y(csr_gpr_iu_rs1_6_) );
	NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__7_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_3503_) );
	MUX2X1 MUX2X1_66 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__7_), .B(csr_gpr_iu_gpr_29__7_), .S(biu_ins_15_bF_buf2), .Y(_3504_) );
	OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .B(_3127__bF_buf0), .C(_3503_), .Y(_3505_) );
	NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf4), .B(_3505_), .Y(_3506_) );
	INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__7_), .Y(_3507_) );
	INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__7_), .Y(_3508_) );
	OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3113__bF_buf6), .C(_3507_), .D(_3105__bF_buf7), .Y(_3509_) );
	INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__7_), .Y(_3510_) );
	INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__7_), .Y(_3511_) );
	OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3110__bF_buf10), .C(_3510_), .D(_3111__bF_buf6), .Y(_3512_) );
	OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3509_), .C(_3117__bF_buf5), .Y(_3513_) );
	NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf7), .B(_3513_), .C(_3506_), .Y(_3514_) );
	NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__7_), .B(_3095__bF_buf2), .Y(_3515_) );
	OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_2811_), .B(_3111__bF_buf5), .C(_3515_), .Y(_3516_) );
	OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_3110__bF_buf9), .C(_2746_), .D(_3113__bF_buf5), .Y(_3517_) );
	OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .B(_3516_), .C(_3109__bF_buf3), .Y(_3518_) );
	INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__7_), .Y(_3519_) );
	INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__7_), .Y(_3520_) );
	OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3111__bF_buf4), .C(_3519_), .D(_3105__bF_buf6), .Y(_3521_) );
	INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__7_), .Y(_3522_) );
	OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3110__bF_buf8), .C(_3522_), .D(_3113__bF_buf4), .Y(_3523_) );
	OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3521_), .C(_3117__bF_buf4), .Y(_3524_) );
	NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_3524_), .B(_3518_), .C(_3107__bF_buf2), .Y(_3525_) );
	NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3525_), .C(_3514_), .Y(_3526_) );
	INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__7_), .Y(_3527_) );
	INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__7_), .Y(_3528_) );
	OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_3111__bF_buf3), .C(_3528_), .D(_3105__bF_buf5), .Y(_3529_) );
	INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__7_), .Y(_3530_) );
	INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__7_), .Y(_3531_) );
	OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3110__bF_buf7), .C(_3530_), .D(_3113__bF_buf3), .Y(_3532_) );
	OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_3529_), .C(_3109__bF_buf2), .Y(_3533_) );
	INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__7_), .Y(_3534_) );
	INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__7_), .Y(_3535_) );
	OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3534_), .B(_3113__bF_buf2), .C(_3535_), .D(_3105__bF_buf4), .Y(_3536_) );
	INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__7_), .Y(_3537_) );
	INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__7_), .Y(_3538_) );
	OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .B(_3110__bF_buf6), .C(_3537_), .D(_3111__bF_buf2), .Y(_3539_) );
	OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_3539_), .B(_3536_), .C(_3117__bF_buf3), .Y(_3540_) );
	AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3533_), .D(_3540_), .Y(_3541_) );
	INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__7_), .Y(_3542_) );
	INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__7_), .Y(_3543_) );
	OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3111__bF_buf1), .C(_3543_), .D(_3105__bF_buf3), .Y(_3544_) );
	INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__7_), .Y(_3545_) );
	INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__7_), .Y(_3546_) );
	OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_3110__bF_buf5), .C(_3545_), .D(_3113__bF_buf1), .Y(_3547_) );
	OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3544_), .C(_3109__bF_buf1), .Y(_3548_) );
	INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__7_), .Y(_3549_) );
	INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__7_), .Y(_3550_) );
	OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_3111__bF_buf0), .C(_3550_), .D(_3105__bF_buf2), .Y(_3551_) );
	INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__7_), .Y(_3552_) );
	INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__7_), .Y(_3553_) );
	OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3110__bF_buf4), .C(_3552_), .D(_3113__bF_buf0), .Y(_3554_) );
	OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_3554_), .B(_3551_), .C(_3117__bF_buf2), .Y(_3555_) );
	AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3548_), .C(_3107__bF_buf1), .Y(_3556_) );
	OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .B(_3556_), .C(_3156__bF_buf2), .Y(_3557_) );
	AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3526_), .D(_3557_), .Y(csr_gpr_iu_rs1_7_) );
	NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__8_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_3558_) );
	MUX2X1 MUX2X1_67 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__8_), .B(csr_gpr_iu_gpr_29__8_), .S(biu_ins_15_bF_buf1), .Y(_3559_) );
	OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3127__bF_buf5), .C(_3558_), .Y(_3560_) );
	NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf0), .B(_3560_), .Y(_3561_) );
	INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__8_), .Y(_3562_) );
	NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__8_), .B(_3095__bF_buf1), .Y(_3563_) );
	OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_3113__bF_buf14), .C(_3563_), .Y(_3564_) );
	INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__8_), .Y(_3565_) );
	INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__8_), .Y(_3566_) );
	OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_3566_), .B(_3110__bF_buf3), .C(_3565_), .D(_3111__bF_buf14), .Y(_3567_) );
	OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_3567_), .B(_3564_), .C(_3117__bF_buf1), .Y(_3568_) );
	NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf6), .B(_3568_), .C(_3561_), .Y(_3569_) );
	NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__8_), .B(_3095__bF_buf0), .Y(_3570_) );
	OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_3111__bF_buf13), .C(_3570_), .Y(_3571_) );
	OAI22X1 OAI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_3110__bF_buf2), .C(_2748_), .D(_3113__bF_buf13), .Y(_3572_) );
	OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3571_), .C(_3109__bF_buf10), .Y(_3573_) );
	INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__8_), .Y(_3574_) );
	NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__8_), .B(_3095__bF_buf11), .Y(_3575_) );
	OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3111__bF_buf12), .C(_3575_), .Y(_3576_) );
	INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__8_), .Y(_3577_) );
	OAI22X1 OAI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3011_), .B(_3110__bF_buf1), .C(_3577_), .D(_3113__bF_buf12), .Y(_3578_) );
	OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(_3576_), .C(_3117__bF_buf0), .Y(_3579_) );
	NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3579_), .C(_3107__bF_buf0), .Y(_3580_) );
	NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3580_), .C(_3569_), .Y(_3581_) );
	INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__8_), .Y(_3582_) );
	INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__8_), .Y(_3583_) );
	OAI22X1 OAI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3110__bF_buf0), .C(_3582_), .D(_3111__bF_buf11), .Y(_3584_) );
	INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__8_), .Y(_3585_) );
	NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__8_), .B(_3095__bF_buf10), .Y(_3586_) );
	OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_3585_), .B(_3113__bF_buf11), .C(_3586_), .Y(_3587_) );
	OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_3584_), .B(_3587_), .C(_3109__bF_buf9), .Y(_3588_) );
	INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__8_), .Y(_3589_) );
	NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__8_), .B(_3095__bF_buf9), .Y(_3590_) );
	OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_3589_), .B(_3113__bF_buf10), .C(_3590_), .Y(_3591_) );
	INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__8_), .Y(_3592_) );
	INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__8_), .Y(_3593_) );
	OAI22X1 OAI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(_3110__bF_buf13), .C(_3592_), .D(_3111__bF_buf10), .Y(_3594_) );
	OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_3594_), .B(_3591_), .C(_3117__bF_buf9), .Y(_3595_) );
	AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3588_), .D(_3595_), .Y(_3596_) );
	INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__8_), .Y(_3597_) );
	INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__8_), .Y(_3598_) );
	OAI22X1 OAI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3110__bF_buf12), .C(_3597_), .D(_3111__bF_buf9), .Y(_3599_) );
	INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__8_), .Y(_3600_) );
	NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__8_), .B(_3095__bF_buf8), .Y(_3601_) );
	OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3113__bF_buf9), .C(_3601_), .Y(_3602_) );
	OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .B(_3602_), .C(_3109__bF_buf8), .Y(_3603_) );
	INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__8_), .Y(_3604_) );
	INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__8_), .Y(_3605_) );
	OAI22X1 OAI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3110__bF_buf11), .C(_3604_), .D(_3111__bF_buf8), .Y(_3606_) );
	INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__8_), .Y(_3607_) );
	NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__8_), .B(_3095__bF_buf7), .Y(_3608_) );
	OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .B(_3113__bF_buf8), .C(_3608_), .Y(_3609_) );
	OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(_3609_), .C(_3117__bF_buf8), .Y(_3610_) );
	AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_3603_), .B(_3610_), .C(_3107__bF_buf5), .Y(_3611_) );
	OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_3596_), .B(_3611_), .C(_3156__bF_buf1), .Y(_3612_) );
	AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3581_), .D(_3612_), .Y(csr_gpr_iu_rs1_8_) );
	NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__9_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_3613_) );
	MUX2X1 MUX2X1_68 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__9_), .B(csr_gpr_iu_gpr_29__9_), .S(biu_ins_15_bF_buf0), .Y(_3614_) );
	OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_3614_), .B(_3127__bF_buf4), .C(_3613_), .Y(_3615_) );
	NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf7), .B(_3615_), .Y(_3616_) );
	INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__9_), .Y(_3617_) );
	NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__9_), .B(_3095__bF_buf6), .Y(_3618_) );
	OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3113__bF_buf6), .C(_3618_), .Y(_3619_) );
	INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__9_), .Y(_3620_) );
	INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__9_), .Y(_3621_) );
	OAI22X1 OAI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3110__bF_buf10), .C(_3620_), .D(_3111__bF_buf6), .Y(_3622_) );
	OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(_3619_), .C(_3117__bF_buf7), .Y(_3623_) );
	NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf5), .B(_3623_), .C(_3616_), .Y(_3624_) );
	NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__9_), .B(_3095__bF_buf5), .Y(_3625_) );
	OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_3111__bF_buf5), .C(_3625_), .Y(_3626_) );
	OAI22X1 OAI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_3110__bF_buf9), .C(_2750_), .D(_3113__bF_buf5), .Y(_3627_) );
	OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_3627_), .B(_3626_), .C(_3109__bF_buf6), .Y(_3628_) );
	INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__9_), .Y(_3629_) );
	NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__9_), .B(_3095__bF_buf4), .Y(_3630_) );
	OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(_3111__bF_buf4), .C(_3630_), .Y(_3631_) );
	INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__9_), .Y(_3632_) );
	OAI22X1 OAI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_3110__bF_buf8), .C(_3632_), .D(_3113__bF_buf4), .Y(_3633_) );
	OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_3633_), .B(_3631_), .C(_3117__bF_buf6), .Y(_3634_) );
	NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_3628_), .B(_3634_), .C(_3107__bF_buf4), .Y(_3635_) );
	NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3635_), .C(_3624_), .Y(_3636_) );
	INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__9_), .Y(_3637_) );
	NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__9_), .B(_3095__bF_buf3), .Y(_3638_) );
	OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3111__bF_buf3), .C(_3638_), .Y(_3639_) );
	INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__9_), .Y(_3640_) );
	INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__9_), .Y(_3641_) );
	OAI22X1 OAI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3110__bF_buf7), .C(_3640_), .D(_3113__bF_buf3), .Y(_3642_) );
	OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3639_), .C(_3109__bF_buf5), .Y(_3643_) );
	INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__9_), .Y(_3644_) );
	INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__9_), .Y(_3645_) );
	OAI22X1 OAI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_3110__bF_buf6), .C(_3644_), .D(_3113__bF_buf2), .Y(_3646_) );
	INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__9_), .Y(_3647_) );
	NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__9_), .B(_3095__bF_buf2), .Y(_3648_) );
	OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3111__bF_buf2), .C(_3648_), .Y(_3649_) );
	OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3649_), .C(_3117__bF_buf5), .Y(_3650_) );
	AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3643_), .D(_3650_), .Y(_3651_) );
	INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__9_), .Y(_3652_) );
	INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__9_), .Y(_3653_) );
	OAI22X1 OAI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3653_), .B(_3110__bF_buf5), .C(_3652_), .D(_3111__bF_buf1), .Y(_3654_) );
	INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__9_), .Y(_3655_) );
	NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__9_), .B(_3095__bF_buf1), .Y(_3656_) );
	OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(_3113__bF_buf1), .C(_3656_), .Y(_3657_) );
	OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_3654_), .B(_3657_), .C(_3109__bF_buf4), .Y(_3658_) );
	INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__9_), .Y(_3659_) );
	INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__9_), .Y(_3660_) );
	OAI22X1 OAI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_3110__bF_buf4), .C(_3659_), .D(_3111__bF_buf0), .Y(_3661_) );
	INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__9_), .Y(_3662_) );
	NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__9_), .B(_3095__bF_buf0), .Y(_3663_) );
	OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_3113__bF_buf0), .C(_3663_), .Y(_3664_) );
	OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3664_), .C(_3117__bF_buf4), .Y(_3665_) );
	AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3665_), .C(_3107__bF_buf3), .Y(_3666_) );
	OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(_3666_), .C(_3156__bF_buf0), .Y(_3667_) );
	AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3636_), .D(_3667_), .Y(csr_gpr_iu_rs1_9_) );
	INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__10_), .Y(_3668_) );
	NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__10_), .B(_3095__bF_buf11), .Y(_3669_) );
	OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .B(_3110__bF_buf3), .C(_3669_), .Y(_3670_) );
	INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__10_), .Y(_3671_) );
	INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__10_), .Y(_3672_) );
	OAI22X1 OAI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3111__bF_buf15), .C(_3672_), .D(_3113__bF_buf15), .Y(_3673_) );
	OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_3673_), .B(_3670_), .C(_3109__bF_buf3), .Y(_3674_) );
	INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__10_), .Y(_3675_) );
	NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__10_), .B(_3095__bF_buf10), .Y(_3676_) );
	OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(_3110__bF_buf2), .C(_3676_), .Y(_3677_) );
	INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__10_), .Y(_3678_) );
	INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__10_), .Y(_3679_) );
	OAI22X1 OAI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3678_), .B(_3111__bF_buf14), .C(_3679_), .D(_3113__bF_buf14), .Y(_3680_) );
	OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_3677_), .C(_3117__bF_buf3), .Y(_3681_) );
	AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3681_), .C(_3107__bF_buf2), .Y(_3682_) );
	INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__10_), .Y(_3683_) );
	INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__10_), .Y(_3684_) );
	OAI22X1 OAI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3111__bF_buf13), .C(_3684_), .D(_3113__bF_buf13), .Y(_3685_) );
	INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__10_), .Y(_3686_) );
	NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__10_), .B(_3095__bF_buf9), .Y(_3687_) );
	OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_3110__bF_buf1), .C(_3687_), .Y(_3688_) );
	OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .B(_3688_), .C(_3109__bF_buf2), .Y(_3689_) );
	INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__10_), .Y(_3690_) );
	INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__10_), .Y(_3691_) );
	OAI22X1 OAI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3690_), .B(_3111__bF_buf12), .C(_3691_), .D(_3113__bF_buf12), .Y(_3692_) );
	INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__10_), .Y(_3693_) );
	NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__10_), .B(_3095__bF_buf8), .Y(_3694_) );
	OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3110__bF_buf0), .C(_3694_), .Y(_3695_) );
	OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .B(_3695_), .C(_3117__bF_buf2), .Y(_3696_) );
	AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_3689_), .B(_3696_), .C(_3126__bF_buf4), .Y(_3697_) );
	OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3697_), .C(_3156__bF_buf4), .Y(_3698_) );
	INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__10_), .Y(_3699_) );
	INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__10_), .Y(_3700_) );
	OAI22X1 OAI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3111__bF_buf11), .C(_3700_), .D(_3113__bF_buf11), .Y(_3701_) );
	AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__10_), .B(_3127__bF_buf3), .C(_3701_), .Y(_3702_) );
	INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__10_), .Y(_3703_) );
	NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__10_), .B(_3095__bF_buf7), .Y(_3704_) );
	OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3113__bF_buf10), .C(_3704_), .Y(_3705_) );
	INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__10_), .Y(_3706_) );
	INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__10_), .Y(_3707_) );
	OAI22X1 OAI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3110__bF_buf13), .C(_3706_), .D(_3111__bF_buf10), .Y(_3708_) );
	OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_3708_), .B(_3705_), .C(_3117__bF_buf1), .Y(_3709_) );
	OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_3117__bF_buf0), .B(_3702_), .C(_3709_), .Y(_3710_) );
	NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__10_), .B(_3095__bF_buf6), .Y(_3711_) );
	OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(_3111__bF_buf9), .C(_3711_), .Y(_3712_) );
	OAI22X1 OAI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_3110__bF_buf12), .C(_2752_), .D(_3113__bF_buf9), .Y(_3713_) );
	OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_3713_), .B(_3712_), .C(_3109__bF_buf1), .Y(_3714_) );
	INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__10_), .Y(_3715_) );
	INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__10_), .Y(_3716_) );
	OAI22X1 OAI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3111__bF_buf8), .C(_3716_), .D(_3113__bF_buf8), .Y(_3717_) );
	NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__10_), .B(_3095__bF_buf5), .Y(_3718_) );
	OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_3015_), .B(_3110__bF_buf11), .C(_3718_), .Y(_3719_) );
	OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .B(_3719_), .C(_3117__bF_buf9), .Y(_3720_) );
	AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_3714_), .B(_3720_), .C(_3126__bF_buf3), .Y(_3721_) );
	AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .B(_3126__bF_buf2), .C(_3721_), .Y(_3722_) );
	OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf2), .B(_3722_), .C(_3698_), .Y(csr_gpr_iu_rs1_10_) );
	INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__11_), .Y(_3723_) );
	NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__11_), .B(_3095__bF_buf4), .Y(_3724_) );
	OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_3110__bF_buf10), .C(_3724_), .Y(_3725_) );
	INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__11_), .Y(_3726_) );
	INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__11_), .Y(_3727_) );
	OAI22X1 OAI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_3111__bF_buf7), .C(_3727_), .D(_3113__bF_buf7), .Y(_3728_) );
	OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_3728_), .B(_3725_), .C(_3109__bF_buf0), .Y(_3729_) );
	INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__11_), .Y(_3730_) );
	NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__11_), .B(_3095__bF_buf3), .Y(_3731_) );
	OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3110__bF_buf9), .C(_3731_), .Y(_3732_) );
	INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__11_), .Y(_3733_) );
	INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__11_), .Y(_3734_) );
	OAI22X1 OAI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3733_), .B(_3111__bF_buf6), .C(_3734_), .D(_3113__bF_buf6), .Y(_3735_) );
	OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .B(_3732_), .C(_3117__bF_buf8), .Y(_3736_) );
	AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .B(_3736_), .C(_3107__bF_buf1), .Y(_3737_) );
	INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__11_), .Y(_3738_) );
	INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__11_), .Y(_3739_) );
	OAI22X1 OAI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3110__bF_buf8), .C(_3738_), .D(_3113__bF_buf5), .Y(_3740_) );
	INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__11_), .Y(_3741_) );
	NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__11_), .B(_3095__bF_buf2), .Y(_3742_) );
	OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_3741_), .B(_3111__bF_buf5), .C(_3742_), .Y(_3743_) );
	OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .B(_3743_), .C(_3109__bF_buf10), .Y(_3744_) );
	INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__11_), .Y(_3745_) );
	INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__11_), .Y(_3746_) );
	OAI22X1 OAI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .B(_3110__bF_buf7), .C(_3745_), .D(_3113__bF_buf4), .Y(_3747_) );
	INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__11_), .Y(_3748_) );
	NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__11_), .B(_3095__bF_buf1), .Y(_3749_) );
	OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3111__bF_buf4), .C(_3749_), .Y(_3750_) );
	OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .B(_3750_), .C(_3117__bF_buf7), .Y(_3751_) );
	AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_3744_), .B(_3751_), .C(_3126__bF_buf1), .Y(_3752_) );
	OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_3737_), .B(_3752_), .C(_3156__bF_buf3), .Y(_3753_) );
	INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__11_), .Y(_3754_) );
	INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__11_), .Y(_3755_) );
	OAI22X1 OAI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3754_), .B(_3111__bF_buf3), .C(_3755_), .D(_3113__bF_buf3), .Y(_3756_) );
	AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__11_), .B(_3127__bF_buf2), .C(_3756_), .Y(_3757_) );
	INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__11_), .Y(_3758_) );
	NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__11_), .B(_3095__bF_buf0), .Y(_3759_) );
	OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_3113__bF_buf2), .C(_3759_), .Y(_3760_) );
	INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__11_), .Y(_3761_) );
	INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__11_), .Y(_3762_) );
	OAI22X1 OAI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_3110__bF_buf6), .C(_3761_), .D(_3111__bF_buf2), .Y(_3763_) );
	OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_3763_), .B(_3760_), .C(_3117__bF_buf6), .Y(_3764_) );
	OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_3117__bF_buf5), .B(_3757_), .C(_3764_), .Y(_3765_) );
	OAI22X1 OAI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_3110__bF_buf5), .C(_2819_), .D(_3111__bF_buf1), .Y(_3766_) );
	NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__11_), .B(_3095__bF_buf11), .Y(_3767_) );
	OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_3113__bF_buf1), .C(_3767_), .Y(_3768_) );
	OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_3766_), .B(_3768_), .C(_3109__bF_buf9), .Y(_3769_) );
	INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__11_), .Y(_3770_) );
	INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__11_), .Y(_3771_) );
	OAI22X1 OAI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3770_), .B(_3111__bF_buf0), .C(_3771_), .D(_3113__bF_buf0), .Y(_3772_) );
	NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__11_), .B(_3095__bF_buf10), .Y(_3773_) );
	OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .B(_3110__bF_buf4), .C(_3773_), .Y(_3774_) );
	OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_3772_), .B(_3774_), .C(_3117__bF_buf4), .Y(_3775_) );
	AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_3769_), .B(_3775_), .C(_3126__bF_buf0), .Y(_3776_) );
	AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(_3126__bF_buf7), .C(_3776_), .Y(_3777_) );
	OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf1), .B(_3777_), .C(_3753_), .Y(csr_gpr_iu_rs1_11_) );
	NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__12_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_3778_) );
	MUX2X1 MUX2X1_69 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__12_), .B(csr_gpr_iu_gpr_29__12_), .S(biu_ins_15_bF_buf6), .Y(_3779_) );
	OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_3127__bF_buf1), .C(_3778_), .Y(_3780_) );
	NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf8), .B(_3780_), .Y(_3781_) );
	INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__12_), .Y(_3782_) );
	NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__12_), .B(_3095__bF_buf9), .Y(_3783_) );
	OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_3113__bF_buf14), .C(_3783_), .Y(_3784_) );
	INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__12_), .Y(_3785_) );
	INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__12_), .Y(_3786_) );
	OAI22X1 OAI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_3110__bF_buf3), .C(_3785_), .D(_3111__bF_buf14), .Y(_3787_) );
	OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(_3784_), .C(_3117__bF_buf3), .Y(_3788_) );
	NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf6), .B(_3788_), .C(_3781_), .Y(_3789_) );
	OAI22X1 OAI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .B(_3110__bF_buf2), .C(_2821_), .D(_3111__bF_buf13), .Y(_3790_) );
	NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__12_), .B(_3095__bF_buf8), .Y(_3791_) );
	OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_3113__bF_buf13), .C(_3791_), .Y(_3792_) );
	OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_3790_), .B(_3792_), .C(_3109__bF_buf7), .Y(_3793_) );
	INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__12_), .Y(_3794_) );
	OAI22X1 OAI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3110__bF_buf1), .C(_3794_), .D(_3111__bF_buf12), .Y(_3795_) );
	INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__12_), .Y(_3796_) );
	NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__12_), .B(_3095__bF_buf7), .Y(_3797_) );
	OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_3113__bF_buf12), .C(_3797_), .Y(_3798_) );
	OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_3798_), .C(_3117__bF_buf2), .Y(_3799_) );
	NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3793_), .B(_3799_), .C(_3107__bF_buf0), .Y(_3800_) );
	NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3800_), .C(_3789_), .Y(_3801_) );
	INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__12_), .Y(_3802_) );
	INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__12_), .Y(_3803_) );
	OAI22X1 OAI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(_3110__bF_buf0), .C(_3802_), .D(_3111__bF_buf11), .Y(_3804_) );
	INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__12_), .Y(_3805_) );
	NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__12_), .B(_3095__bF_buf6), .Y(_3806_) );
	OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3113__bF_buf11), .C(_3806_), .Y(_3807_) );
	OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(_3807_), .C(_3109__bF_buf6), .Y(_3808_) );
	INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__12_), .Y(_3809_) );
	NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__12_), .B(_3095__bF_buf5), .Y(_3810_) );
	OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_3809_), .B(_3113__bF_buf10), .C(_3810_), .Y(_3811_) );
	INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__12_), .Y(_3812_) );
	INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__12_), .Y(_3813_) );
	OAI22X1 OAI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_3110__bF_buf13), .C(_3812_), .D(_3111__bF_buf10), .Y(_3814_) );
	OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_3814_), .B(_3811_), .C(_3117__bF_buf1), .Y(_3815_) );
	AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_3808_), .D(_3815_), .Y(_3816_) );
	INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__12_), .Y(_3817_) );
	NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__12_), .B(_3095__bF_buf4), .Y(_3818_) );
	OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(_3111__bF_buf9), .C(_3818_), .Y(_3819_) );
	INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__12_), .Y(_3820_) );
	INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__12_), .Y(_3821_) );
	OAI22X1 OAI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_3110__bF_buf12), .C(_3820_), .D(_3113__bF_buf9), .Y(_3822_) );
	OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_3822_), .B(_3819_), .C(_3109__bF_buf5), .Y(_3823_) );
	INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__12_), .Y(_3824_) );
	NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__12_), .B(_3095__bF_buf3), .Y(_3825_) );
	OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_3111__bF_buf8), .C(_3825_), .Y(_3826_) );
	INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__12_), .Y(_3827_) );
	INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__12_), .Y(_3828_) );
	OAI22X1 OAI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_3110__bF_buf11), .C(_3827_), .D(_3113__bF_buf8), .Y(_3829_) );
	OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3826_), .C(_3117__bF_buf0), .Y(_3830_) );
	AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_3823_), .B(_3830_), .C(_3107__bF_buf5), .Y(_3831_) );
	OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .B(_3831_), .C(_3156__bF_buf2), .Y(_3832_) );
	AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_3801_), .D(_3832_), .Y(csr_gpr_iu_rs1_12_) );
	INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__13_), .Y(_3833_) );
	INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__13_), .Y(_3834_) );
	OAI22X1 OAI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(_3110__bF_buf10), .C(_3833_), .D(_3105__bF_buf1), .Y(_3835_) );
	INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__13_), .Y(_3836_) );
	INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__13_), .Y(_3837_) );
	OAI22X1 OAI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_3111__bF_buf7), .C(_3837_), .D(_3113__bF_buf7), .Y(_3838_) );
	OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3838_), .C(_3109__bF_buf4), .Y(_3839_) );
	INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__13_), .Y(_3840_) );
	INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__13_), .Y(_3841_) );
	OAI22X1 OAI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3110__bF_buf9), .C(_3840_), .D(_3105__bF_buf0), .Y(_3842_) );
	INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__13_), .Y(_3843_) );
	INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__13_), .Y(_3844_) );
	OAI22X1 OAI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_3111__bF_buf6), .C(_3844_), .D(_3113__bF_buf6), .Y(_3845_) );
	OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_3842_), .B(_3845_), .C(_3117__bF_buf9), .Y(_3846_) );
	AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3839_), .C(_3107__bF_buf4), .Y(_3847_) );
	INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__13_), .Y(_3848_) );
	NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__13_), .B(_3095__bF_buf2), .Y(_3849_) );
	OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .B(_3113__bF_buf5), .C(_3849_), .Y(_3850_) );
	INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__13_), .Y(_3851_) );
	INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__13_), .Y(_3852_) );
	OAI22X1 OAI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_3110__bF_buf8), .C(_3851_), .D(_3111__bF_buf5), .Y(_3853_) );
	OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3850_), .C(_3109__bF_buf3), .Y(_3854_) );
	INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__13_), .Y(_3855_) );
	NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__13_), .B(_3095__bF_buf1), .Y(_3856_) );
	OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .B(_3113__bF_buf4), .C(_3856_), .Y(_3857_) );
	INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__13_), .Y(_3858_) );
	INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__13_), .Y(_3859_) );
	OAI22X1 OAI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(_3110__bF_buf7), .C(_3858_), .D(_3111__bF_buf4), .Y(_3860_) );
	OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .B(_3857_), .C(_3117__bF_buf8), .Y(_3861_) );
	AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_3854_), .B(_3861_), .C(_3126__bF_buf5), .Y(_3862_) );
	OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(_3862_), .C(_3156__bF_buf1), .Y(_3863_) );
	INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__13_), .Y(_3864_) );
	INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__13_), .Y(_3865_) );
	OAI22X1 OAI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .B(_3111__bF_buf3), .C(_3865_), .D(_3113__bF_buf3), .Y(_3866_) );
	INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__13_), .Y(_3867_) );
	NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__13_), .B(biu_ins_15_bF_buf5), .Y(_3868_) );
	OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf4), .B(_3867_), .C(_3868_), .Y(_3869_) );
	AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf0), .B(_3869_), .C(_3866_), .Y(_3870_) );
	INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__13_), .Y(_3871_) );
	INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__13_), .Y(_3872_) );
	OAI22X1 OAI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3111__bF_buf2), .C(_3872_), .D(_3113__bF_buf2), .Y(_3873_) );
	AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__13_), .B(_3127__bF_buf5), .C(_3873_), .Y(_3874_) );
	MUX2X1 MUX2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3874_), .B(_3870_), .S(_3109__bF_buf2), .Y(_3875_) );
	NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__13_), .B(_3095__bF_buf0), .Y(_3876_) );
	OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_3111__bF_buf1), .C(_3876_), .Y(_3877_) );
	OAI22X1 OAI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_3110__bF_buf6), .C(_2758_), .D(_3113__bF_buf1), .Y(_3878_) );
	OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_3878_), .B(_3877_), .C(_3109__bF_buf1), .Y(_3879_) );
	INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__13_), .Y(_3880_) );
	INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__13_), .Y(_3881_) );
	OAI22X1 OAI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_3880_), .B(_3111__bF_buf0), .C(_3881_), .D(_3113__bF_buf0), .Y(_3882_) );
	INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__13_), .Y(_3883_) );
	OAI22X1 OAI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3110__bF_buf5), .C(_3883_), .D(_3105__bF_buf7), .Y(_3884_) );
	OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_3884_), .B(_3882_), .C(_3117__bF_buf7), .Y(_3885_) );
	AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_3879_), .B(_3885_), .C(_3126__bF_buf4), .Y(_3886_) );
	AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .B(_3126__bF_buf3), .C(_3886_), .Y(_3887_) );
	OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf0), .B(_3887_), .C(_3863_), .Y(csr_gpr_iu_rs1_13_) );
	INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__14_), .Y(_3888_) );
	INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__14_), .Y(_3889_) );
	OAI22X1 OAI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_3110__bF_buf4), .C(_3888_), .D(_3105__bF_buf6), .Y(_3890_) );
	INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__14_), .Y(_3891_) );
	INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__14_), .Y(_3892_) );
	OAI22X1 OAI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_3111__bF_buf15), .C(_3892_), .D(_3113__bF_buf15), .Y(_3893_) );
	OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_3890_), .B(_3893_), .C(_3109__bF_buf0), .Y(_3894_) );
	INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__14_), .Y(_3895_) );
	INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__14_), .Y(_3896_) );
	OAI22X1 OAI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_3896_), .B(_3110__bF_buf3), .C(_3895_), .D(_3105__bF_buf5), .Y(_3897_) );
	INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__14_), .Y(_3898_) );
	INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__14_), .Y(_3899_) );
	OAI22X1 OAI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(_3111__bF_buf14), .C(_3899_), .D(_3113__bF_buf14), .Y(_3900_) );
	OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3900_), .C(_3117__bF_buf6), .Y(_3901_) );
	AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_3894_), .C(_3107__bF_buf3), .Y(_3902_) );
	INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__14_), .Y(_3903_) );
	INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__14_), .Y(_3904_) );
	OAI22X1 OAI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3904_), .B(_3110__bF_buf2), .C(_3903_), .D(_3113__bF_buf13), .Y(_3905_) );
	INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__14_), .Y(_3906_) );
	NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__14_), .B(_3095__bF_buf11), .Y(_3907_) );
	OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3111__bF_buf13), .C(_3907_), .Y(_3908_) );
	OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_3905_), .B(_3908_), .C(_3109__bF_buf10), .Y(_3909_) );
	INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__14_), .Y(_3910_) );
	INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__14_), .Y(_3911_) );
	OAI22X1 OAI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_3110__bF_buf1), .C(_3910_), .D(_3113__bF_buf12), .Y(_3912_) );
	INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__14_), .Y(_3913_) );
	NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__14_), .B(_3095__bF_buf10), .Y(_3914_) );
	OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3111__bF_buf12), .C(_3914_), .Y(_3915_) );
	OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3915_), .C(_3117__bF_buf5), .Y(_3916_) );
	AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_3909_), .B(_3916_), .C(_3126__bF_buf2), .Y(_3917_) );
	OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .B(_3917_), .C(_3156__bF_buf0), .Y(_3918_) );
	INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__14_), .Y(_3919_) );
	INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__14_), .Y(_3920_) );
	OAI22X1 OAI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_3111__bF_buf11), .C(_3920_), .D(_3113__bF_buf11), .Y(_3921_) );
	INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__14_), .Y(_3922_) );
	NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__14_), .B(biu_ins_15_bF_buf3), .Y(_3923_) );
	OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf2), .B(_3922_), .C(_3923_), .Y(_3924_) );
	AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf4), .B(_3924_), .C(_3921_), .Y(_3925_) );
	INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__14_), .Y(_3926_) );
	INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__14_), .Y(_3927_) );
	OAI22X1 OAI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_3111__bF_buf10), .C(_3927_), .D(_3113__bF_buf10), .Y(_3928_) );
	AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__14_), .B(_3127__bF_buf3), .C(_3928_), .Y(_3929_) );
	MUX2X1 MUX2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3929_), .B(_3925_), .S(_3109__bF_buf9), .Y(_3930_) );
	OAI22X1 OAI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_3110__bF_buf0), .C(_2825_), .D(_3111__bF_buf9), .Y(_3931_) );
	NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__14_), .B(_3095__bF_buf9), .Y(_3932_) );
	OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_3113__bF_buf9), .C(_3932_), .Y(_3933_) );
	OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_3931_), .B(_3933_), .C(_3109__bF_buf8), .Y(_3934_) );
	INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__14_), .Y(_3935_) );
	INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__14_), .Y(_3936_) );
	OAI22X1 OAI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3111__bF_buf8), .C(_3936_), .D(_3113__bF_buf8), .Y(_3937_) );
	INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__14_), .Y(_3938_) );
	OAI22X1 OAI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_3110__bF_buf13), .C(_3938_), .D(_3105__bF_buf4), .Y(_3939_) );
	OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_3939_), .B(_3937_), .C(_3117__bF_buf4), .Y(_3940_) );
	AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_3934_), .B(_3940_), .C(_3126__bF_buf1), .Y(_3941_) );
	AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_3126__bF_buf0), .C(_3941_), .Y(_3942_) );
	OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf3), .B(_3942_), .C(_3918_), .Y(csr_gpr_iu_rs1_14_) );
	INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__15_), .Y(_3943_) );
	INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__15_), .Y(_3944_) );
	OAI22X1 OAI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3944_), .B(_3110__bF_buf12), .C(_3943_), .D(_3105__bF_buf3), .Y(_3945_) );
	INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__15_), .Y(_3946_) );
	INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__15_), .Y(_3947_) );
	OAI22X1 OAI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_3111__bF_buf7), .C(_3947_), .D(_3113__bF_buf7), .Y(_3948_) );
	OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_3945_), .B(_3948_), .C(_3109__bF_buf7), .Y(_3949_) );
	INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__15_), .Y(_3950_) );
	INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__15_), .Y(_3951_) );
	OAI22X1 OAI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3110__bF_buf11), .C(_3950_), .D(_3105__bF_buf2), .Y(_3952_) );
	INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__15_), .Y(_3953_) );
	INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__15_), .Y(_3954_) );
	OAI22X1 OAI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_3111__bF_buf6), .C(_3954_), .D(_3113__bF_buf6), .Y(_3955_) );
	OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .B(_3955_), .C(_3117__bF_buf3), .Y(_3956_) );
	AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_3949_), .C(_3107__bF_buf2), .Y(_3957_) );
	INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__15_), .Y(_3958_) );
	INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__15_), .Y(_3959_) );
	OAI22X1 OAI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_3110__bF_buf10), .C(_3958_), .D(_3113__bF_buf5), .Y(_3960_) );
	INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__15_), .Y(_3961_) );
	NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__15_), .B(_3095__bF_buf8), .Y(_3962_) );
	OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_3111__bF_buf5), .C(_3962_), .Y(_3963_) );
	OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_3960_), .B(_3963_), .C(_3109__bF_buf6), .Y(_3964_) );
	INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__15_), .Y(_3965_) );
	INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__15_), .Y(_3966_) );
	OAI22X1 OAI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(_3966_), .B(_3110__bF_buf9), .C(_3965_), .D(_3113__bF_buf4), .Y(_3967_) );
	INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__15_), .Y(_3968_) );
	NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__15_), .B(_3095__bF_buf7), .Y(_3969_) );
	OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3111__bF_buf4), .C(_3969_), .Y(_3970_) );
	OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_3970_), .C(_3117__bF_buf2), .Y(_3971_) );
	AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .B(_3971_), .C(_3126__bF_buf7), .Y(_3972_) );
	OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_3957_), .B(_3972_), .C(_3156__bF_buf4), .Y(_3973_) );
	INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__15_), .Y(_3974_) );
	INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__15_), .Y(_3975_) );
	OAI22X1 OAI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_3974_), .B(_3111__bF_buf3), .C(_3975_), .D(_3113__bF_buf3), .Y(_3976_) );
	INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__15_), .Y(_3977_) );
	NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__15_), .B(biu_ins_15_bF_buf1), .Y(_3978_) );
	OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf0), .B(_3977_), .C(_3978_), .Y(_3979_) );
	AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf2), .B(_3979_), .C(_3976_), .Y(_3980_) );
	INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__15_), .Y(_3981_) );
	INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__15_), .Y(_3982_) );
	OAI22X1 OAI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(_3981_), .B(_3111__bF_buf2), .C(_3982_), .D(_3113__bF_buf2), .Y(_3983_) );
	AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__15_), .B(_3127__bF_buf1), .C(_3983_), .Y(_3984_) );
	MUX2X1 MUX2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3984_), .B(_3980_), .S(_3109__bF_buf5), .Y(_3985_) );
	NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__15_), .B(_3095__bF_buf6), .Y(_3986_) );
	OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_3111__bF_buf1), .C(_3986_), .Y(_3987_) );
	OAI22X1 OAI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_2892_), .B(_3110__bF_buf8), .C(_2762_), .D(_3113__bF_buf1), .Y(_3988_) );
	OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(_3987_), .C(_3109__bF_buf4), .Y(_3989_) );
	INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__15_), .Y(_3990_) );
	INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__15_), .Y(_3991_) );
	OAI22X1 OAI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_3111__bF_buf0), .C(_3991_), .D(_3113__bF_buf0), .Y(_3992_) );
	INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__15_), .Y(_3993_) );
	OAI22X1 OAI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3110__bF_buf7), .C(_3993_), .D(_3105__bF_buf1), .Y(_3994_) );
	OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_3994_), .B(_3992_), .C(_3117__bF_buf1), .Y(_3995_) );
	AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_3995_), .C(_3126__bF_buf6), .Y(_3996_) );
	AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_3985_), .B(_3126__bF_buf5), .C(_3996_), .Y(_3997_) );
	OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf2), .B(_3997_), .C(_3973_), .Y(csr_gpr_iu_rs1_15_) );
	NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__16_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_3998_) );
	MUX2X1 MUX2X1_73 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__16_), .B(csr_gpr_iu_gpr_29__16_), .S(biu_ins_15_bF_buf6), .Y(_3999_) );
	OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_3999_), .B(_3127__bF_buf0), .C(_3998_), .Y(_4000_) );
	NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf3), .B(_4000_), .Y(_4001_) );
	INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__16_), .Y(_4002_) );
	NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__16_), .B(_3095__bF_buf5), .Y(_4003_) );
	OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_4002_), .B(_3113__bF_buf14), .C(_4003_), .Y(_4004_) );
	INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__16_), .Y(_4005_) );
	INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__16_), .Y(_4006_) );
	OAI22X1 OAI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_3110__bF_buf6), .C(_4005_), .D(_3111__bF_buf14), .Y(_4007_) );
	OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_4007_), .B(_4004_), .C(_3117__bF_buf0), .Y(_4008_) );
	NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf4), .B(_4008_), .C(_4001_), .Y(_4009_) );
	OAI22X1 OAI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_3110__bF_buf5), .C(_2829_), .D(_3111__bF_buf13), .Y(_4010_) );
	NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__16_), .B(_3095__bF_buf4), .Y(_4011_) );
	OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_2764_), .B(_3113__bF_buf13), .C(_4011_), .Y(_4012_) );
	OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4012_), .C(_3109__bF_buf2), .Y(_4013_) );
	INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__16_), .Y(_4014_) );
	OAI22X1 OAI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_3110__bF_buf4), .C(_4014_), .D(_3111__bF_buf12), .Y(_4015_) );
	INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__16_), .Y(_4016_) );
	NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__16_), .B(_3095__bF_buf3), .Y(_4017_) );
	OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_4016_), .B(_3113__bF_buf12), .C(_4017_), .Y(_4018_) );
	OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_4015_), .B(_4018_), .C(_3117__bF_buf9), .Y(_4019_) );
	NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_4013_), .B(_4019_), .C(_3107__bF_buf1), .Y(_4020_) );
	NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4020_), .C(_4009_), .Y(_4021_) );
	INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__16_), .Y(_4022_) );
	NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__16_), .B(_3095__bF_buf2), .Y(_4023_) );
	OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_3111__bF_buf11), .C(_4023_), .Y(_4024_) );
	INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__16_), .Y(_4025_) );
	INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__16_), .Y(_4026_) );
	OAI22X1 OAI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .B(_3110__bF_buf3), .C(_4025_), .D(_3113__bF_buf11), .Y(_4027_) );
	OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(_4024_), .C(_3109__bF_buf1), .Y(_4028_) );
	INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__16_), .Y(_4029_) );
	NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__16_), .B(_3095__bF_buf1), .Y(_4030_) );
	OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_4029_), .B(_3113__bF_buf10), .C(_4030_), .Y(_4031_) );
	INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__16_), .Y(_4032_) );
	INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__16_), .Y(_4033_) );
	OAI22X1 OAI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .B(_3110__bF_buf2), .C(_4032_), .D(_3111__bF_buf10), .Y(_4034_) );
	OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .B(_4031_), .C(_3117__bF_buf8), .Y(_4035_) );
	AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4028_), .D(_4035_), .Y(_4036_) );
	INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__16_), .Y(_4037_) );
	NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__16_), .B(_3095__bF_buf0), .Y(_4038_) );
	OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(_3111__bF_buf9), .C(_4038_), .Y(_4039_) );
	INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__16_), .Y(_4040_) );
	INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__16_), .Y(_4041_) );
	OAI22X1 OAI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(_4041_), .B(_3110__bF_buf1), .C(_4040_), .D(_3113__bF_buf9), .Y(_4042_) );
	OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4039_), .C(_3109__bF_buf0), .Y(_4043_) );
	INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__16_), .Y(_4044_) );
	NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__16_), .B(_3095__bF_buf11), .Y(_4045_) );
	OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_4044_), .B(_3111__bF_buf8), .C(_4045_), .Y(_4046_) );
	INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__16_), .Y(_4047_) );
	INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__16_), .Y(_4048_) );
	OAI22X1 OAI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_3110__bF_buf0), .C(_4047_), .D(_3113__bF_buf8), .Y(_4049_) );
	OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_4049_), .B(_4046_), .C(_3117__bF_buf7), .Y(_4050_) );
	AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4043_), .B(_4050_), .C(_3107__bF_buf0), .Y(_4051_) );
	OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .B(_4051_), .C(_3156__bF_buf3), .Y(_4052_) );
	AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4021_), .D(_4052_), .Y(csr_gpr_iu_rs1_16_) );
	NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__17_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_4053_) );
	MUX2X1 MUX2X1_74 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__17_), .B(csr_gpr_iu_gpr_29__17_), .S(biu_ins_15_bF_buf5), .Y(_4054_) );
	OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_3127__bF_buf5), .C(_4053_), .Y(_4055_) );
	NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf10), .B(_4055_), .Y(_4056_) );
	INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__17_), .Y(_4057_) );
	NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__17_), .B(_3095__bF_buf10), .Y(_4058_) );
	OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .B(_3113__bF_buf6), .C(_4058_), .Y(_4059_) );
	INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__17_), .Y(_4060_) );
	INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__17_), .Y(_4061_) );
	OAI22X1 OAI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(_4061_), .B(_3110__bF_buf13), .C(_4060_), .D(_3111__bF_buf6), .Y(_4062_) );
	OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_4062_), .B(_4059_), .C(_3117__bF_buf6), .Y(_4063_) );
	NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf3), .B(_4063_), .C(_4056_), .Y(_4064_) );
	NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__17_), .B(_3095__bF_buf9), .Y(_4065_) );
	OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_3111__bF_buf5), .C(_4065_), .Y(_4066_) );
	OAI22X1 OAI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_3110__bF_buf12), .C(_2766_), .D(_3113__bF_buf5), .Y(_4067_) );
	OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_4067_), .B(_4066_), .C(_3109__bF_buf9), .Y(_4068_) );
	INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__17_), .Y(_4069_) );
	NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__17_), .B(_3095__bF_buf8), .Y(_4070_) );
	OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_3111__bF_buf4), .C(_4070_), .Y(_4071_) );
	INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__17_), .Y(_4072_) );
	OAI22X1 OAI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .B(_3110__bF_buf11), .C(_4072_), .D(_3113__bF_buf4), .Y(_4073_) );
	OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(_4071_), .C(_3117__bF_buf5), .Y(_4074_) );
	NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_4074_), .C(_3107__bF_buf5), .Y(_4075_) );
	NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4075_), .C(_4064_), .Y(_4076_) );
	INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__17_), .Y(_4077_) );
	NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__17_), .B(_3095__bF_buf7), .Y(_4078_) );
	OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_4077_), .B(_3111__bF_buf3), .C(_4078_), .Y(_4079_) );
	INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__17_), .Y(_4080_) );
	INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__17_), .Y(_4081_) );
	OAI22X1 OAI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(_3110__bF_buf10), .C(_4080_), .D(_3113__bF_buf3), .Y(_4082_) );
	OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_4082_), .B(_4079_), .C(_3109__bF_buf8), .Y(_4083_) );
	INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__17_), .Y(_4084_) );
	NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__17_), .B(_3095__bF_buf6), .Y(_4085_) );
	OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .B(_3113__bF_buf2), .C(_4085_), .Y(_4086_) );
	INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__17_), .Y(_4087_) );
	INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__17_), .Y(_4088_) );
	OAI22X1 OAI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .B(_3110__bF_buf9), .C(_4087_), .D(_3111__bF_buf2), .Y(_4089_) );
	OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_4089_), .B(_4086_), .C(_3117__bF_buf4), .Y(_4090_) );
	AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4083_), .D(_4090_), .Y(_4091_) );
	INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__17_), .Y(_4092_) );
	NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__17_), .B(_3095__bF_buf5), .Y(_4093_) );
	OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_4092_), .B(_3111__bF_buf1), .C(_4093_), .Y(_4094_) );
	INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__17_), .Y(_4095_) );
	INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__17_), .Y(_4096_) );
	OAI22X1 OAI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_3110__bF_buf8), .C(_4095_), .D(_3113__bF_buf1), .Y(_4097_) );
	OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_4097_), .B(_4094_), .C(_3109__bF_buf7), .Y(_4098_) );
	INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__17_), .Y(_4099_) );
	NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__17_), .B(_3095__bF_buf4), .Y(_4100_) );
	OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_3111__bF_buf0), .C(_4100_), .Y(_4101_) );
	INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__17_), .Y(_4102_) );
	INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__17_), .Y(_4103_) );
	OAI22X1 OAI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .B(_3110__bF_buf7), .C(_4102_), .D(_3113__bF_buf0), .Y(_4104_) );
	OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_4104_), .B(_4101_), .C(_3117__bF_buf3), .Y(_4105_) );
	AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_4098_), .B(_4105_), .C(_3107__bF_buf4), .Y(_4106_) );
	OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_4091_), .B(_4106_), .C(_3156__bF_buf2), .Y(_4107_) );
	AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4076_), .D(_4107_), .Y(csr_gpr_iu_rs1_17_) );
	NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__18_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_4108_) );
	MUX2X1 MUX2X1_75 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__18_), .B(csr_gpr_iu_gpr_29__18_), .S(biu_ins_15_bF_buf4), .Y(_4109_) );
	OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_4109_), .B(_3127__bF_buf4), .C(_4108_), .Y(_4110_) );
	NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf6), .B(_4110_), .Y(_4111_) );
	INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__18_), .Y(_4112_) );
	INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__18_), .Y(_4113_) );
	OAI22X1 OAI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .B(_3113__bF_buf14), .C(_4112_), .D(_3105__bF_buf0), .Y(_4114_) );
	INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__18_), .Y(_4115_) );
	INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__18_), .Y(_4116_) );
	OAI22X1 OAI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .B(_3110__bF_buf6), .C(_4115_), .D(_3111__bF_buf14), .Y(_4117_) );
	OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .B(_4114_), .C(_3117__bF_buf2), .Y(_4118_) );
	NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf2), .B(_4118_), .C(_4111_), .Y(_4119_) );
	OAI22X1 OAI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_3110__bF_buf5), .C(_2833_), .D(_3111__bF_buf13), .Y(_4120_) );
	NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__18_), .B(_3095__bF_buf3), .Y(_4121_) );
	OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_3113__bF_buf13), .C(_4121_), .Y(_4122_) );
	OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_4120_), .B(_4122_), .C(_3109__bF_buf5), .Y(_4123_) );
	INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__18_), .Y(_4124_) );
	OAI22X1 OAI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_3110__bF_buf4), .C(_4124_), .D(_3111__bF_buf12), .Y(_4125_) );
	INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__18_), .Y(_4126_) );
	INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__18_), .Y(_4127_) );
	OAI22X1 OAI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(_4127_), .B(_3113__bF_buf12), .C(_4126_), .D(_3105__bF_buf7), .Y(_4128_) );
	OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_4125_), .B(_4128_), .C(_3117__bF_buf1), .Y(_4129_) );
	NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_4129_), .B(_4123_), .C(_3107__bF_buf3), .Y(_4130_) );
	NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4130_), .C(_4119_), .Y(_4131_) );
	INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__18_), .Y(_4132_) );
	NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__18_), .B(_3095__bF_buf2), .Y(_4133_) );
	OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_4132_), .B(_3111__bF_buf11), .C(_4133_), .Y(_4134_) );
	INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__18_), .Y(_4135_) );
	INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__18_), .Y(_4136_) );
	OAI22X1 OAI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_3110__bF_buf3), .C(_4135_), .D(_3113__bF_buf11), .Y(_4137_) );
	OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_4137_), .B(_4134_), .C(_3109__bF_buf4), .Y(_4138_) );
	INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__18_), .Y(_4139_) );
	NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__18_), .B(_3095__bF_buf1), .Y(_4140_) );
	OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_3113__bF_buf10), .C(_4140_), .Y(_4141_) );
	INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__18_), .Y(_4142_) );
	INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__18_), .Y(_4143_) );
	OAI22X1 OAI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(_4143_), .B(_3110__bF_buf2), .C(_4142_), .D(_3111__bF_buf10), .Y(_4144_) );
	OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(_4141_), .C(_3117__bF_buf0), .Y(_4145_) );
	AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4138_), .D(_4145_), .Y(_4146_) );
	INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__18_), .Y(_4147_) );
	INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__18_), .Y(_4148_) );
	OAI22X1 OAI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_3110__bF_buf1), .C(_4147_), .D(_3111__bF_buf9), .Y(_4149_) );
	INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__18_), .Y(_4150_) );
	INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__18_), .Y(_4151_) );
	OAI22X1 OAI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(_4150_), .B(_3113__bF_buf9), .C(_4151_), .D(_3105__bF_buf6), .Y(_4152_) );
	OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_4149_), .B(_4152_), .C(_3109__bF_buf3), .Y(_4153_) );
	INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__18_), .Y(_4154_) );
	INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__18_), .Y(_4155_) );
	OAI22X1 OAI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_3110__bF_buf0), .C(_4154_), .D(_3111__bF_buf8), .Y(_4156_) );
	INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__18_), .Y(_4157_) );
	INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__18_), .Y(_4158_) );
	OAI22X1 OAI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(_4157_), .B(_3113__bF_buf8), .C(_4158_), .D(_3105__bF_buf5), .Y(_4159_) );
	OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_4156_), .B(_4159_), .C(_3117__bF_buf9), .Y(_4160_) );
	AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_4153_), .C(_3107__bF_buf2), .Y(_4161_) );
	OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4161_), .C(_3156__bF_buf1), .Y(_4162_) );
	AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4131_), .D(_4162_), .Y(csr_gpr_iu_rs1_18_) );
	INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__19_), .Y(_4163_) );
	INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__19_), .Y(_4164_) );
	OAI22X1 OAI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(_4164_), .B(_3110__bF_buf13), .C(_4163_), .D(_3105__bF_buf4), .Y(_4165_) );
	INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__19_), .Y(_4166_) );
	INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__19_), .Y(_4167_) );
	OAI22X1 OAI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_3111__bF_buf7), .C(_4167_), .D(_3113__bF_buf7), .Y(_4168_) );
	OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4168_), .C(_3109__bF_buf2), .Y(_4169_) );
	INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__19_), .Y(_4170_) );
	INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__19_), .Y(_4171_) );
	OAI22X1 OAI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .B(_3110__bF_buf12), .C(_4170_), .D(_3105__bF_buf3), .Y(_4172_) );
	INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__19_), .Y(_4173_) );
	INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__19_), .Y(_4174_) );
	OAI22X1 OAI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_3111__bF_buf6), .C(_4174_), .D(_3113__bF_buf6), .Y(_4175_) );
	OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4175_), .C(_3117__bF_buf8), .Y(_4176_) );
	AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_4176_), .B(_4169_), .C(_3107__bF_buf1), .Y(_4177_) );
	INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__19_), .Y(_4178_) );
	NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__19_), .B(_3095__bF_buf0), .Y(_4179_) );
	OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_3113__bF_buf5), .C(_4179_), .Y(_4180_) );
	INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__19_), .Y(_4181_) );
	INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__19_), .Y(_4182_) );
	OAI22X1 OAI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .B(_3110__bF_buf11), .C(_4181_), .D(_3111__bF_buf5), .Y(_4183_) );
	OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_4183_), .B(_4180_), .C(_3109__bF_buf1), .Y(_4184_) );
	INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__19_), .Y(_4185_) );
	NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__19_), .B(_3095__bF_buf11), .Y(_4186_) );
	OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_4185_), .B(_3113__bF_buf4), .C(_4186_), .Y(_4187_) );
	INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__19_), .Y(_4188_) );
	INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__19_), .Y(_4189_) );
	OAI22X1 OAI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .B(_3110__bF_buf10), .C(_4188_), .D(_3111__bF_buf4), .Y(_4190_) );
	OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_4190_), .B(_4187_), .C(_3117__bF_buf7), .Y(_4191_) );
	AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4184_), .B(_4191_), .C(_3126__bF_buf1), .Y(_4192_) );
	OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_4177_), .B(_4192_), .C(_3156__bF_buf0), .Y(_4193_) );
	INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__19_), .Y(_4194_) );
	INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__19_), .Y(_4195_) );
	OAI22X1 OAI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(_4194_), .B(_3111__bF_buf3), .C(_4195_), .D(_3113__bF_buf3), .Y(_4196_) );
	INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__19_), .Y(_4197_) );
	NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__19_), .B(biu_ins_15_bF_buf3), .Y(_4198_) );
	OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf2), .B(_4197_), .C(_4198_), .Y(_4199_) );
	AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf3), .B(_4199_), .C(_4196_), .Y(_4200_) );
	INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__19_), .Y(_4201_) );
	INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__19_), .Y(_4202_) );
	OAI22X1 OAI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(_4201_), .B(_3111__bF_buf2), .C(_4202_), .D(_3113__bF_buf2), .Y(_4203_) );
	AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__19_), .B(_3127__bF_buf2), .C(_4203_), .Y(_4204_) );
	MUX2X1 MUX2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_4204_), .B(_4200_), .S(_3109__bF_buf0), .Y(_4205_) );
	NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__19_), .B(_3095__bF_buf10), .Y(_4206_) );
	OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .B(_3111__bF_buf1), .C(_4206_), .Y(_4207_) );
	OAI22X1 OAI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_3110__bF_buf9), .C(_2770_), .D(_3113__bF_buf1), .Y(_4208_) );
	OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_4208_), .B(_4207_), .C(_3109__bF_buf10), .Y(_4209_) );
	INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__19_), .Y(_4210_) );
	INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__19_), .Y(_4211_) );
	OAI22X1 OAI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(_4210_), .B(_3111__bF_buf0), .C(_4211_), .D(_3113__bF_buf0), .Y(_4212_) );
	INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__19_), .Y(_4213_) );
	OAI22X1 OAI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .B(_3110__bF_buf8), .C(_4213_), .D(_3105__bF_buf2), .Y(_4214_) );
	OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_4214_), .B(_4212_), .C(_3117__bF_buf6), .Y(_4215_) );
	AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_4209_), .B(_4215_), .C(_3126__bF_buf0), .Y(_4216_) );
	AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_4205_), .B(_3126__bF_buf7), .C(_4216_), .Y(_4217_) );
	OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf1), .B(_4217_), .C(_4193_), .Y(csr_gpr_iu_rs1_19_) );
	NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__20_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_4218_) );
	MUX2X1 MUX2X1_77 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__20_), .B(csr_gpr_iu_gpr_29__20_), .S(biu_ins_15_bF_buf1), .Y(_4219_) );
	OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_4219_), .B(_3127__bF_buf1), .C(_4218_), .Y(_4220_) );
	NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf9), .B(_4220_), .Y(_4221_) );
	INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__20_), .Y(_4222_) );
	NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__20_), .B(_3095__bF_buf9), .Y(_4223_) );
	OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_4222_), .B(_3113__bF_buf14), .C(_4223_), .Y(_4224_) );
	INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__20_), .Y(_4225_) );
	INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__20_), .Y(_4226_) );
	OAI22X1 OAI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_3110__bF_buf7), .C(_4225_), .D(_3111__bF_buf14), .Y(_4227_) );
	OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_4227_), .B(_4224_), .C(_3117__bF_buf5), .Y(_4228_) );
	NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf6), .B(_4228_), .C(_4221_), .Y(_4229_) );
	OAI22X1 OAI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_3110__bF_buf6), .C(_2837_), .D(_3111__bF_buf13), .Y(_4230_) );
	NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__20_), .B(_3095__bF_buf8), .Y(_4231_) );
	OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_3113__bF_buf13), .C(_4231_), .Y(_4232_) );
	OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_4230_), .B(_4232_), .C(_3109__bF_buf8), .Y(_4233_) );
	INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__20_), .Y(_4234_) );
	OAI22X1 OAI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_3110__bF_buf5), .C(_4234_), .D(_3111__bF_buf12), .Y(_4235_) );
	INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__20_), .Y(_4236_) );
	NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__20_), .B(_3095__bF_buf7), .Y(_4237_) );
	OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_3113__bF_buf12), .C(_4237_), .Y(_4238_) );
	OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_4235_), .B(_4238_), .C(_3117__bF_buf4), .Y(_4239_) );
	NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_4233_), .B(_4239_), .C(_3107__bF_buf0), .Y(_4240_) );
	NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4240_), .C(_4229_), .Y(_4241_) );
	INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__20_), .Y(_4242_) );
	NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__20_), .B(_3095__bF_buf6), .Y(_4243_) );
	OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_4242_), .B(_3111__bF_buf11), .C(_4243_), .Y(_4244_) );
	INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__20_), .Y(_4245_) );
	INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__20_), .Y(_4246_) );
	OAI22X1 OAI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(_4246_), .B(_3110__bF_buf4), .C(_4245_), .D(_3113__bF_buf11), .Y(_4247_) );
	OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_4247_), .B(_4244_), .C(_3109__bF_buf7), .Y(_4248_) );
	INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__20_), .Y(_4249_) );
	INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__20_), .Y(_4250_) );
	OAI22X1 OAI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(_4250_), .B(_3110__bF_buf3), .C(_4249_), .D(_3113__bF_buf10), .Y(_4251_) );
	INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__20_), .Y(_4252_) );
	NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__20_), .B(_3095__bF_buf5), .Y(_4253_) );
	OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_4252_), .B(_3111__bF_buf10), .C(_4253_), .Y(_4254_) );
	OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_4251_), .B(_4254_), .C(_3117__bF_buf3), .Y(_4255_) );
	AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4248_), .D(_4255_), .Y(_4256_) );
	INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__20_), .Y(_4257_) );
	NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__20_), .B(_3095__bF_buf4), .Y(_4258_) );
	OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_4257_), .B(_3111__bF_buf9), .C(_4258_), .Y(_4259_) );
	INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__20_), .Y(_4260_) );
	INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__20_), .Y(_4261_) );
	OAI22X1 OAI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(_3110__bF_buf2), .C(_4260_), .D(_3113__bF_buf9), .Y(_4262_) );
	OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_4262_), .B(_4259_), .C(_3109__bF_buf6), .Y(_4263_) );
	INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__20_), .Y(_4264_) );
	NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__20_), .B(_3095__bF_buf3), .Y(_4265_) );
	OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_4264_), .B(_3111__bF_buf8), .C(_4265_), .Y(_4266_) );
	INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__20_), .Y(_4267_) );
	INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__20_), .Y(_4268_) );
	OAI22X1 OAI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(_4268_), .B(_3110__bF_buf1), .C(_4267_), .D(_3113__bF_buf8), .Y(_4269_) );
	OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .B(_4266_), .C(_3117__bF_buf2), .Y(_4270_) );
	AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_4263_), .B(_4270_), .C(_3107__bF_buf5), .Y(_4271_) );
	OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_4256_), .B(_4271_), .C(_3156__bF_buf4), .Y(_4272_) );
	AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4241_), .D(_4272_), .Y(csr_gpr_iu_rs1_20_) );
	INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__21_), .Y(_4273_) );
	INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__21_), .Y(_4274_) );
	OAI22X1 OAI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(_4274_), .B(_3110__bF_buf0), .C(_4273_), .D(_3105__bF_buf1), .Y(_4275_) );
	INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__21_), .Y(_4276_) );
	INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__21_), .Y(_4277_) );
	OAI22X1 OAI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(_4276_), .B(_3111__bF_buf7), .C(_4277_), .D(_3113__bF_buf7), .Y(_4278_) );
	OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_4275_), .B(_4278_), .C(_3109__bF_buf5), .Y(_4279_) );
	INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__21_), .Y(_4280_) );
	INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__21_), .Y(_4281_) );
	OAI22X1 OAI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_3110__bF_buf13), .C(_4280_), .D(_3105__bF_buf0), .Y(_4282_) );
	INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__21_), .Y(_4283_) );
	INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__21_), .Y(_4284_) );
	OAI22X1 OAI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(_4283_), .B(_3111__bF_buf6), .C(_4284_), .D(_3113__bF_buf6), .Y(_4285_) );
	OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_4282_), .B(_4285_), .C(_3117__bF_buf1), .Y(_4286_) );
	AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(_4279_), .C(_3107__bF_buf4), .Y(_4287_) );
	INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__21_), .Y(_4288_) );
	INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__21_), .Y(_4289_) );
	OAI22X1 OAI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(_4288_), .B(_3111__bF_buf5), .C(_4289_), .D(_3113__bF_buf5), .Y(_4290_) );
	INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__21_), .Y(_4291_) );
	INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__21_), .Y(_4292_) );
	OAI22X1 OAI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .B(_3110__bF_buf12), .C(_4291_), .D(_3105__bF_buf7), .Y(_4293_) );
	OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(_4290_), .C(_3109__bF_buf4), .Y(_4294_) );
	INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__21_), .Y(_4295_) );
	INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__21_), .Y(_4296_) );
	OAI22X1 OAI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(_4295_), .B(_3111__bF_buf4), .C(_4296_), .D(_3113__bF_buf4), .Y(_4297_) );
	INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__21_), .Y(_4298_) );
	INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__21_), .Y(_4299_) );
	OAI22X1 OAI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(_4299_), .B(_3110__bF_buf11), .C(_4298_), .D(_3105__bF_buf6), .Y(_4300_) );
	OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_4300_), .B(_4297_), .C(_3117__bF_buf0), .Y(_4301_) );
	AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_4301_), .B(_4294_), .C(_3126__bF_buf5), .Y(_4302_) );
	OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_4302_), .C(_3156__bF_buf3), .Y(_4303_) );
	INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__21_), .Y(_4304_) );
	INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__21_), .Y(_4305_) );
	OAI22X1 OAI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(_4304_), .B(_3111__bF_buf3), .C(_4305_), .D(_3113__bF_buf3), .Y(_4306_) );
	INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__21_), .Y(_4307_) );
	NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__21_), .B(biu_ins_15_bF_buf0), .Y(_4308_) );
	OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf6), .B(_4307_), .C(_4308_), .Y(_4309_) );
	AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf0), .B(_4309_), .C(_4306_), .Y(_4310_) );
	INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__21_), .Y(_4311_) );
	INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__21_), .Y(_4312_) );
	OAI22X1 OAI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(_4311_), .B(_3111__bF_buf2), .C(_4312_), .D(_3113__bF_buf2), .Y(_4313_) );
	AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__21_), .B(_3127__bF_buf5), .C(_4313_), .Y(_4314_) );
	MUX2X1 MUX2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_4310_), .S(_3109__bF_buf3), .Y(_4315_) );
	OAI22X1 OAI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(_3110__bF_buf10), .C(_2839_), .D(_3111__bF_buf1), .Y(_4316_) );
	NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__21_), .B(_3095__bF_buf2), .Y(_4317_) );
	OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .B(_3113__bF_buf1), .C(_4317_), .Y(_4318_) );
	OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_4316_), .B(_4318_), .C(_3109__bF_buf2), .Y(_4319_) );
	INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__21_), .Y(_4320_) );
	INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__21_), .Y(_4321_) );
	OAI22X1 OAI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(_4320_), .B(_3111__bF_buf0), .C(_4321_), .D(_3113__bF_buf0), .Y(_4322_) );
	INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__21_), .Y(_4323_) );
	OAI22X1 OAI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_3110__bF_buf9), .C(_4323_), .D(_3105__bF_buf5), .Y(_4324_) );
	OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_4324_), .B(_4322_), .C(_3117__bF_buf9), .Y(_4325_) );
	AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_4319_), .B(_4325_), .C(_3126__bF_buf4), .Y(_4326_) );
	AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .B(_3126__bF_buf3), .C(_4326_), .Y(_4327_) );
	OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf0), .B(_4327_), .C(_4303_), .Y(csr_gpr_iu_rs1_21_) );
	INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__22_), .Y(_4328_) );
	NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__22_), .B(_3095__bF_buf1), .Y(_4329_) );
	OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_4328_), .B(_3110__bF_buf8), .C(_4329_), .Y(_4330_) );
	INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__22_), .Y(_4331_) );
	INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__22_), .Y(_4332_) );
	OAI22X1 OAI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(_3111__bF_buf15), .C(_4332_), .D(_3113__bF_buf15), .Y(_4333_) );
	OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_4333_), .B(_4330_), .C(_3109__bF_buf1), .Y(_4334_) );
	INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__22_), .Y(_4335_) );
	NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__22_), .B(_3095__bF_buf0), .Y(_4336_) );
	OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_3110__bF_buf7), .C(_4336_), .Y(_4337_) );
	INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__22_), .Y(_4338_) );
	INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__22_), .Y(_4339_) );
	OAI22X1 OAI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(_4338_), .B(_3111__bF_buf14), .C(_4339_), .D(_3113__bF_buf14), .Y(_4340_) );
	OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4337_), .C(_3117__bF_buf8), .Y(_4341_) );
	AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4334_), .B(_4341_), .C(_3107__bF_buf3), .Y(_4342_) );
	INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__22_), .Y(_4343_) );
	NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__22_), .B(_3095__bF_buf11), .Y(_4344_) );
	OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_3113__bF_buf13), .C(_4344_), .Y(_4345_) );
	INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__22_), .Y(_4346_) );
	INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__22_), .Y(_4347_) );
	OAI22X1 OAI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .B(_3110__bF_buf6), .C(_4346_), .D(_3111__bF_buf13), .Y(_4348_) );
	OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_4348_), .B(_4345_), .C(_3109__bF_buf0), .Y(_4349_) );
	INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__22_), .Y(_4350_) );
	NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__22_), .B(_3095__bF_buf10), .Y(_4351_) );
	OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_3113__bF_buf12), .C(_4351_), .Y(_4352_) );
	INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__22_), .Y(_4353_) );
	INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__22_), .Y(_4354_) );
	OAI22X1 OAI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_3110__bF_buf5), .C(_4353_), .D(_3111__bF_buf12), .Y(_4355_) );
	OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_4355_), .B(_4352_), .C(_3117__bF_buf7), .Y(_4356_) );
	AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_4349_), .B(_4356_), .C(_3126__bF_buf2), .Y(_4357_) );
	OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_4342_), .B(_4357_), .C(_3156__bF_buf2), .Y(_4358_) );
	INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__22_), .Y(_4359_) );
	INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__22_), .Y(_4360_) );
	OAI22X1 OAI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(_4359_), .B(_3111__bF_buf11), .C(_4360_), .D(_3113__bF_buf11), .Y(_4361_) );
	AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__22_), .B(_3127__bF_buf4), .C(_4361_), .Y(_4362_) );
	INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__22_), .Y(_4363_) );
	NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__22_), .B(_3095__bF_buf9), .Y(_4364_) );
	OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_4363_), .B(_3113__bF_buf10), .C(_4364_), .Y(_4365_) );
	INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__22_), .Y(_4366_) );
	INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__22_), .Y(_4367_) );
	OAI22X1 OAI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(_4367_), .B(_3110__bF_buf4), .C(_4366_), .D(_3111__bF_buf10), .Y(_4368_) );
	OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_4368_), .B(_4365_), .C(_3117__bF_buf6), .Y(_4369_) );
	OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_3117__bF_buf5), .B(_4362_), .C(_4369_), .Y(_4370_) );
	NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__22_), .B(_3095__bF_buf8), .Y(_4371_) );
	OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_2841_), .B(_3111__bF_buf9), .C(_4371_), .Y(_4372_) );
	OAI22X1 OAI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .B(_3110__bF_buf3), .C(_2776_), .D(_3113__bF_buf9), .Y(_4373_) );
	OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_4373_), .B(_4372_), .C(_3109__bF_buf10), .Y(_4374_) );
	INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__22_), .Y(_4375_) );
	INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__22_), .Y(_4376_) );
	OAI22X1 OAI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(_4375_), .B(_3111__bF_buf8), .C(_4376_), .D(_3113__bF_buf8), .Y(_4377_) );
	NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__22_), .B(_3095__bF_buf7), .Y(_4378_) );
	OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .B(_3110__bF_buf2), .C(_4378_), .Y(_4379_) );
	OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_4377_), .B(_4379_), .C(_3117__bF_buf4), .Y(_4380_) );
	AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_4374_), .B(_4380_), .C(_3126__bF_buf1), .Y(_4381_) );
	AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4370_), .B(_3126__bF_buf0), .C(_4381_), .Y(_4382_) );
	OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf3), .B(_4382_), .C(_4358_), .Y(csr_gpr_iu_rs1_22_) );
	INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__23_), .Y(_4383_) );
	INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__23_), .Y(_4384_) );
	OAI22X1 OAI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(_3110__bF_buf1), .C(_4383_), .D(_3105__bF_buf4), .Y(_4385_) );
	INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__23_), .Y(_4386_) );
	INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__23_), .Y(_4387_) );
	OAI22X1 OAI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(_4386_), .B(_3111__bF_buf7), .C(_4387_), .D(_3113__bF_buf7), .Y(_4388_) );
	OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_4388_), .C(_3109__bF_buf9), .Y(_4389_) );
	INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__23_), .Y(_4390_) );
	INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__23_), .Y(_4391_) );
	OAI22X1 OAI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(_4391_), .B(_3110__bF_buf0), .C(_4390_), .D(_3105__bF_buf3), .Y(_4392_) );
	INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__23_), .Y(_4393_) );
	INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__23_), .Y(_4394_) );
	OAI22X1 OAI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3111__bF_buf6), .C(_4394_), .D(_3113__bF_buf6), .Y(_4395_) );
	OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_4392_), .B(_4395_), .C(_3117__bF_buf3), .Y(_4396_) );
	AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_4396_), .B(_4389_), .C(_3107__bF_buf2), .Y(_4397_) );
	INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__23_), .Y(_4398_) );
	INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__23_), .Y(_4399_) );
	OAI22X1 OAI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(_4399_), .B(_3110__bF_buf13), .C(_4398_), .D(_3113__bF_buf5), .Y(_4400_) );
	INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__23_), .Y(_4401_) );
	INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__23_), .Y(_4402_) );
	OAI22X1 OAI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_3111__bF_buf5), .C(_4402_), .D(_3105__bF_buf2), .Y(_4403_) );
	OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_4400_), .B(_4403_), .C(_3109__bF_buf8), .Y(_4404_) );
	INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__23_), .Y(_4405_) );
	INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__23_), .Y(_4406_) );
	OAI22X1 OAI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_3110__bF_buf12), .C(_4405_), .D(_3113__bF_buf4), .Y(_4407_) );
	INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__23_), .Y(_4408_) );
	INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__23_), .Y(_4409_) );
	OAI22X1 OAI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(_4408_), .B(_3111__bF_buf4), .C(_4409_), .D(_3105__bF_buf1), .Y(_4410_) );
	OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_4407_), .B(_4410_), .C(_3117__bF_buf2), .Y(_4411_) );
	AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4411_), .B(_4404_), .C(_3126__bF_buf7), .Y(_4412_) );
	OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_4397_), .B(_4412_), .C(_3156__bF_buf1), .Y(_4413_) );
	INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__23_), .Y(_4414_) );
	INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__23_), .Y(_4415_) );
	OAI22X1 OAI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_3111__bF_buf3), .C(_4415_), .D(_3113__bF_buf3), .Y(_4416_) );
	INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__23_), .Y(_4417_) );
	NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__23_), .B(biu_ins_15_bF_buf5), .Y(_4418_) );
	OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf4), .B(_4417_), .C(_4418_), .Y(_4419_) );
	AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf3), .B(_4419_), .C(_4416_), .Y(_4420_) );
	INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__23_), .Y(_4421_) );
	INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__23_), .Y(_4422_) );
	OAI22X1 OAI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .B(_3111__bF_buf2), .C(_4422_), .D(_3113__bF_buf2), .Y(_4423_) );
	AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__23_), .B(_3127__bF_buf2), .C(_4423_), .Y(_4424_) );
	MUX2X1 MUX2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .B(_4420_), .S(_3109__bF_buf7), .Y(_4425_) );
	OAI22X1 OAI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_3110__bF_buf11), .C(_2843_), .D(_3111__bF_buf1), .Y(_4426_) );
	NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__23_), .B(_3095__bF_buf6), .Y(_4427_) );
	OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_2778_), .B(_3113__bF_buf1), .C(_4427_), .Y(_4428_) );
	OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_4426_), .B(_4428_), .C(_3109__bF_buf6), .Y(_4429_) );
	INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__23_), .Y(_4430_) );
	INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__23_), .Y(_4431_) );
	OAI22X1 OAI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_3111__bF_buf0), .C(_4431_), .D(_3113__bF_buf0), .Y(_4432_) );
	INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__23_), .Y(_4433_) );
	OAI22X1 OAI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3110__bF_buf10), .C(_4433_), .D(_3105__bF_buf0), .Y(_4434_) );
	OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4432_), .C(_3117__bF_buf1), .Y(_4435_) );
	AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4435_), .C(_3126__bF_buf6), .Y(_4436_) );
	AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .B(_3126__bF_buf5), .C(_4436_), .Y(_4437_) );
	OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf2), .B(_4437_), .C(_4413_), .Y(csr_gpr_iu_rs1_23_) );
	NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__24_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_4438_) );
	MUX2X1 MUX2X1_80 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__24_), .B(csr_gpr_iu_gpr_29__24_), .S(biu_ins_15_bF_buf3), .Y(_4439_) );
	OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_4439_), .B(_3127__bF_buf1), .C(_4438_), .Y(_4440_) );
	NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf5), .B(_4440_), .Y(_4441_) );
	INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__24_), .Y(_4442_) );
	NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__24_), .B(_3095__bF_buf5), .Y(_4443_) );
	OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_3113__bF_buf14), .C(_4443_), .Y(_4444_) );
	INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__24_), .Y(_4445_) );
	INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__24_), .Y(_4446_) );
	OAI22X1 OAI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_3110__bF_buf9), .C(_4445_), .D(_3111__bF_buf14), .Y(_4447_) );
	OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_4447_), .B(_4444_), .C(_3117__bF_buf0), .Y(_4448_) );
	NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf4), .B(_4448_), .C(_4441_), .Y(_4449_) );
	OAI22X1 OAI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2910_), .B(_3110__bF_buf8), .C(_2845_), .D(_3111__bF_buf13), .Y(_4450_) );
	NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__24_), .B(_3095__bF_buf4), .Y(_4451_) );
	OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_3113__bF_buf13), .C(_4451_), .Y(_4452_) );
	OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_4450_), .B(_4452_), .C(_3109__bF_buf4), .Y(_4453_) );
	INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__24_), .Y(_4454_) );
	OAI22X1 OAI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_3110__bF_buf7), .C(_4454_), .D(_3111__bF_buf12), .Y(_4455_) );
	INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__24_), .Y(_4456_) );
	NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__24_), .B(_3095__bF_buf3), .Y(_4457_) );
	OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_3113__bF_buf12), .C(_4457_), .Y(_4458_) );
	OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_4455_), .B(_4458_), .C(_3117__bF_buf9), .Y(_4459_) );
	NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_4453_), .B(_4459_), .C(_3107__bF_buf1), .Y(_4460_) );
	NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4460_), .C(_4449_), .Y(_4461_) );
	INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__24_), .Y(_4462_) );
	NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__24_), .B(_3095__bF_buf2), .Y(_4463_) );
	OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_4462_), .B(_3111__bF_buf11), .C(_4463_), .Y(_4464_) );
	INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__24_), .Y(_4465_) );
	INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__24_), .Y(_4466_) );
	OAI22X1 OAI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(_4466_), .B(_3110__bF_buf6), .C(_4465_), .D(_3113__bF_buf11), .Y(_4467_) );
	OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_4467_), .B(_4464_), .C(_3109__bF_buf3), .Y(_4468_) );
	INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__24_), .Y(_4469_) );
	NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__24_), .B(_3095__bF_buf1), .Y(_4470_) );
	OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_4469_), .B(_3113__bF_buf10), .C(_4470_), .Y(_4471_) );
	INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__24_), .Y(_4472_) );
	INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__24_), .Y(_4473_) );
	OAI22X1 OAI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(_4473_), .B(_3110__bF_buf5), .C(_4472_), .D(_3111__bF_buf10), .Y(_4474_) );
	OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_4474_), .B(_4471_), .C(_3117__bF_buf8), .Y(_4475_) );
	AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4468_), .D(_4475_), .Y(_4476_) );
	INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__24_), .Y(_4477_) );
	INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__24_), .Y(_4478_) );
	OAI22X1 OAI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_3110__bF_buf4), .C(_4477_), .D(_3111__bF_buf9), .Y(_4479_) );
	INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__24_), .Y(_4480_) );
	NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__24_), .B(_3095__bF_buf0), .Y(_4481_) );
	OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_3113__bF_buf9), .C(_4481_), .Y(_4482_) );
	OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_4482_), .C(_3109__bF_buf2), .Y(_4483_) );
	INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__24_), .Y(_4484_) );
	INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__24_), .Y(_4485_) );
	OAI22X1 OAI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_3110__bF_buf3), .C(_4484_), .D(_3111__bF_buf8), .Y(_4486_) );
	INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__24_), .Y(_4487_) );
	NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__24_), .B(_3095__bF_buf11), .Y(_4488_) );
	OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_3113__bF_buf8), .C(_4488_), .Y(_4489_) );
	OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_4486_), .B(_4489_), .C(_3117__bF_buf7), .Y(_4490_) );
	AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .B(_4490_), .C(_3107__bF_buf0), .Y(_4491_) );
	OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_4476_), .B(_4491_), .C(_3156__bF_buf0), .Y(_4492_) );
	AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4461_), .D(_4492_), .Y(csr_gpr_iu_rs1_24_) );
	NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__25_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_4493_) );
	MUX2X1 MUX2X1_81 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__25_), .B(csr_gpr_iu_gpr_29__25_), .S(biu_ins_15_bF_buf2), .Y(_4494_) );
	OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_4494_), .B(_3127__bF_buf0), .C(_4493_), .Y(_4495_) );
	NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf1), .B(_4495_), .Y(_4496_) );
	INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__25_), .Y(_4497_) );
	NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__25_), .B(_3095__bF_buf10), .Y(_4498_) );
	OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_4497_), .B(_3113__bF_buf6), .C(_4498_), .Y(_4499_) );
	INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__25_), .Y(_4500_) );
	INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__25_), .Y(_4501_) );
	OAI22X1 OAI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_3110__bF_buf2), .C(_4500_), .D(_3111__bF_buf6), .Y(_4502_) );
	OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_4502_), .B(_4499_), .C(_3117__bF_buf6), .Y(_4503_) );
	NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf3), .B(_4503_), .C(_4496_), .Y(_4504_) );
	NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__25_), .B(_3095__bF_buf9), .Y(_4505_) );
	OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_3111__bF_buf5), .C(_4505_), .Y(_4506_) );
	OAI22X1 OAI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_3110__bF_buf1), .C(_2782_), .D(_3113__bF_buf5), .Y(_4507_) );
	OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_4507_), .B(_4506_), .C(_3109__bF_buf0), .Y(_4508_) );
	INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__25_), .Y(_4509_) );
	NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__25_), .B(_3095__bF_buf8), .Y(_4510_) );
	OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_4509_), .B(_3111__bF_buf4), .C(_4510_), .Y(_4511_) );
	INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__25_), .Y(_4512_) );
	OAI22X1 OAI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3045_), .B(_3110__bF_buf0), .C(_4512_), .D(_3113__bF_buf4), .Y(_4513_) );
	OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_4513_), .B(_4511_), .C(_3117__bF_buf5), .Y(_4514_) );
	NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_4508_), .B(_4514_), .C(_3107__bF_buf5), .Y(_4515_) );
	NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4515_), .C(_4504_), .Y(_4516_) );
	INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__25_), .Y(_4517_) );
	NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__25_), .B(_3095__bF_buf7), .Y(_4518_) );
	OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_4517_), .B(_3111__bF_buf3), .C(_4518_), .Y(_4519_) );
	INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__25_), .Y(_4520_) );
	INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__25_), .Y(_4521_) );
	OAI22X1 OAI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(_4521_), .B(_3110__bF_buf13), .C(_4520_), .D(_3113__bF_buf3), .Y(_4522_) );
	OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_4522_), .B(_4519_), .C(_3109__bF_buf10), .Y(_4523_) );
	INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__25_), .Y(_4524_) );
	NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__25_), .B(_3095__bF_buf6), .Y(_4525_) );
	OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_4524_), .B(_3113__bF_buf2), .C(_4525_), .Y(_4526_) );
	INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__25_), .Y(_4527_) );
	INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__25_), .Y(_4528_) );
	OAI22X1 OAI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(_4528_), .B(_3110__bF_buf12), .C(_4527_), .D(_3111__bF_buf2), .Y(_4529_) );
	OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_4529_), .B(_4526_), .C(_3117__bF_buf4), .Y(_4530_) );
	AOI22X1 AOI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4523_), .D(_4530_), .Y(_4531_) );
	INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__25_), .Y(_4532_) );
	NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__25_), .B(_3095__bF_buf5), .Y(_4533_) );
	OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_4532_), .B(_3111__bF_buf1), .C(_4533_), .Y(_4534_) );
	INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__25_), .Y(_4535_) );
	INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__25_), .Y(_4536_) );
	OAI22X1 OAI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_3110__bF_buf11), .C(_4535_), .D(_3113__bF_buf1), .Y(_4537_) );
	OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_4537_), .B(_4534_), .C(_3109__bF_buf9), .Y(_4538_) );
	INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__25_), .Y(_4539_) );
	NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__25_), .B(_3095__bF_buf4), .Y(_4540_) );
	OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_3111__bF_buf0), .C(_4540_), .Y(_4541_) );
	INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__25_), .Y(_4542_) );
	INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__25_), .Y(_4543_) );
	OAI22X1 OAI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(_4543_), .B(_3110__bF_buf10), .C(_4542_), .D(_3113__bF_buf0), .Y(_4544_) );
	OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_4544_), .B(_4541_), .C(_3117__bF_buf3), .Y(_4545_) );
	AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .B(_4545_), .C(_3107__bF_buf4), .Y(_4546_) );
	OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_4531_), .B(_4546_), .C(_3156__bF_buf4), .Y(_4547_) );
	AOI22X1 AOI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4516_), .D(_4547_), .Y(csr_gpr_iu_rs1_25_) );
	INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__26_), .Y(_4548_) );
	INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__26_), .Y(_4549_) );
	OAI22X1 OAI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(_4549_), .B(_3110__bF_buf9), .C(_4548_), .D(_3105__bF_buf7), .Y(_4550_) );
	INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__26_), .Y(_4551_) );
	INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__26_), .Y(_4552_) );
	OAI22X1 OAI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_3111__bF_buf15), .C(_4552_), .D(_3113__bF_buf15), .Y(_4553_) );
	OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_4550_), .B(_4553_), .C(_3109__bF_buf8), .Y(_4554_) );
	INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__26_), .Y(_4555_) );
	INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__26_), .Y(_4556_) );
	OAI22X1 OAI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_3110__bF_buf8), .C(_4555_), .D(_3105__bF_buf6), .Y(_4557_) );
	INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__26_), .Y(_4558_) );
	INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__26_), .Y(_4559_) );
	OAI22X1 OAI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(_4558_), .B(_3111__bF_buf14), .C(_4559_), .D(_3113__bF_buf14), .Y(_4560_) );
	OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_4557_), .B(_4560_), .C(_3117__bF_buf2), .Y(_4561_) );
	AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_4561_), .B(_4554_), .C(_3107__bF_buf3), .Y(_4562_) );
	INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__26_), .Y(_4563_) );
	INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__26_), .Y(_4564_) );
	OAI22X1 OAI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(_4564_), .B(_3110__bF_buf7), .C(_4563_), .D(_3113__bF_buf13), .Y(_4565_) );
	INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__26_), .Y(_4566_) );
	INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__26_), .Y(_4567_) );
	OAI22X1 OAI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(_4566_), .B(_3111__bF_buf13), .C(_4567_), .D(_3105__bF_buf5), .Y(_4568_) );
	OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_4565_), .B(_4568_), .C(_3109__bF_buf7), .Y(_4569_) );
	INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__26_), .Y(_4570_) );
	INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__26_), .Y(_4571_) );
	OAI22X1 OAI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(_4571_), .B(_3110__bF_buf6), .C(_4570_), .D(_3113__bF_buf12), .Y(_4572_) );
	INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__26_), .Y(_4573_) );
	INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__26_), .Y(_4574_) );
	OAI22X1 OAI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_3111__bF_buf12), .C(_4574_), .D(_3105__bF_buf4), .Y(_4575_) );
	OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_4572_), .B(_4575_), .C(_3117__bF_buf1), .Y(_4576_) );
	AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4569_), .C(_3126__bF_buf2), .Y(_4577_) );
	OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_4577_), .C(_3156__bF_buf3), .Y(_4578_) );
	INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__26_), .Y(_4579_) );
	INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__26_), .Y(_4580_) );
	OAI22X1 OAI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(_4579_), .B(_3111__bF_buf11), .C(_4580_), .D(_3113__bF_buf11), .Y(_4581_) );
	INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__26_), .Y(_4582_) );
	NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__26_), .B(biu_ins_15_bF_buf1), .Y(_4583_) );
	OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf0), .B(_4582_), .C(_4583_), .Y(_4584_) );
	AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf5), .B(_4584_), .C(_4581_), .Y(_4585_) );
	INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__26_), .Y(_4586_) );
	INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__26_), .Y(_4587_) );
	OAI22X1 OAI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_3111__bF_buf10), .C(_4587_), .D(_3113__bF_buf10), .Y(_4588_) );
	AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__26_), .B(_3127__bF_buf4), .C(_4588_), .Y(_4589_) );
	MUX2X1 MUX2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .B(_4585_), .S(_3109__bF_buf6), .Y(_4590_) );
	NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__26_), .B(_3095__bF_buf3), .Y(_4591_) );
	OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_3111__bF_buf9), .C(_4591_), .Y(_4592_) );
	OAI22X1 OAI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_3110__bF_buf5), .C(_2784_), .D(_3113__bF_buf9), .Y(_4593_) );
	OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_4593_), .B(_4592_), .C(_3109__bF_buf5), .Y(_4594_) );
	INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__26_), .Y(_4595_) );
	INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__26_), .Y(_4596_) );
	OAI22X1 OAI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_3111__bF_buf8), .C(_4596_), .D(_3113__bF_buf8), .Y(_4597_) );
	INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__26_), .Y(_4598_) );
	OAI22X1 OAI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_3110__bF_buf4), .C(_4598_), .D(_3105__bF_buf3), .Y(_4599_) );
	OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(_4597_), .C(_3117__bF_buf0), .Y(_4600_) );
	AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .B(_4600_), .C(_3126__bF_buf1), .Y(_4601_) );
	AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_4590_), .B(_3126__bF_buf0), .C(_4601_), .Y(_4602_) );
	OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf1), .B(_4602_), .C(_4578_), .Y(csr_gpr_iu_rs1_26_) );
	INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__27_), .Y(_4603_) );
	INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__27_), .Y(_4604_) );
	OAI22X1 OAI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .B(_3110__bF_buf3), .C(_4603_), .D(_3105__bF_buf2), .Y(_4605_) );
	INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__27_), .Y(_4606_) );
	INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__27_), .Y(_4607_) );
	OAI22X1 OAI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_3111__bF_buf7), .C(_4607_), .D(_3113__bF_buf7), .Y(_4608_) );
	OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_4605_), .B(_4608_), .C(_3109__bF_buf4), .Y(_4609_) );
	INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__27_), .Y(_4610_) );
	INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__27_), .Y(_4611_) );
	OAI22X1 OAI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_3110__bF_buf2), .C(_4610_), .D(_3105__bF_buf1), .Y(_4612_) );
	INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__27_), .Y(_4613_) );
	INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__27_), .Y(_4614_) );
	OAI22X1 OAI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_3111__bF_buf6), .C(_4614_), .D(_3113__bF_buf6), .Y(_4615_) );
	OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_4612_), .B(_4615_), .C(_3117__bF_buf9), .Y(_4616_) );
	AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_4616_), .B(_4609_), .C(_3107__bF_buf2), .Y(_4617_) );
	INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__27_), .Y(_4618_) );
	INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__27_), .Y(_4619_) );
	OAI22X1 OAI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(_4618_), .B(_3111__bF_buf5), .C(_4619_), .D(_3113__bF_buf5), .Y(_4620_) );
	INVX1 INVX1_1005 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__27_), .Y(_4621_) );
	NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__27_), .B(_3095__bF_buf2), .Y(_4622_) );
	OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_3110__bF_buf1), .C(_4622_), .Y(_4623_) );
	OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4623_), .C(_3109__bF_buf3), .Y(_4624_) );
	INVX1 INVX1_1006 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__27_), .Y(_4625_) );
	INVX1 INVX1_1007 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__27_), .Y(_4626_) );
	OAI22X1 OAI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(_4625_), .B(_3111__bF_buf4), .C(_4626_), .D(_3113__bF_buf4), .Y(_4627_) );
	INVX1 INVX1_1008 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__27_), .Y(_4628_) );
	NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__27_), .B(_3095__bF_buf1), .Y(_4629_) );
	OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_3110__bF_buf0), .C(_4629_), .Y(_4630_) );
	OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_4627_), .B(_4630_), .C(_3117__bF_buf8), .Y(_4631_) );
	AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_4624_), .B(_4631_), .C(_3126__bF_buf7), .Y(_4632_) );
	OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4632_), .C(_3156__bF_buf2), .Y(_4633_) );
	INVX1 INVX1_1009 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__27_), .Y(_4634_) );
	INVX1 INVX1_1010 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__27_), .Y(_4635_) );
	OAI22X1 OAI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_3111__bF_buf3), .C(_4635_), .D(_3113__bF_buf3), .Y(_4636_) );
	INVX1 INVX1_1011 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__27_), .Y(_4637_) );
	NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__27_), .B(biu_ins_15_bF_buf6), .Y(_4638_) );
	OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf5), .B(_4637_), .C(_4638_), .Y(_4639_) );
	AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf3), .B(_4639_), .C(_4636_), .Y(_4640_) );
	INVX1 INVX1_1012 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__27_), .Y(_4641_) );
	INVX1 INVX1_1013 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__27_), .Y(_4642_) );
	OAI22X1 OAI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .B(_3111__bF_buf2), .C(_4642_), .D(_3113__bF_buf2), .Y(_4643_) );
	AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__27_), .B(_3127__bF_buf2), .C(_4643_), .Y(_4644_) );
	MUX2X1 MUX2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4644_), .B(_4640_), .S(_3109__bF_buf2), .Y(_4645_) );
	NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__27_), .B(_3095__bF_buf0), .Y(_4646_) );
	OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_2851_), .B(_3111__bF_buf1), .C(_4646_), .Y(_4647_) );
	OAI22X1 OAI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .B(_3110__bF_buf13), .C(_2786_), .D(_3113__bF_buf1), .Y(_4648_) );
	OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_4648_), .B(_4647_), .C(_3109__bF_buf1), .Y(_4649_) );
	INVX1 INVX1_1014 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__27_), .Y(_4650_) );
	INVX1 INVX1_1015 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__27_), .Y(_4651_) );
	OAI22X1 OAI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(_4650_), .B(_3111__bF_buf0), .C(_4651_), .D(_3113__bF_buf0), .Y(_4652_) );
	INVX1 INVX1_1016 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__27_), .Y(_4653_) );
	OAI22X1 OAI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_3110__bF_buf12), .C(_4653_), .D(_3105__bF_buf0), .Y(_4654_) );
	OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4652_), .C(_3117__bF_buf7), .Y(_4655_) );
	AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_4649_), .B(_4655_), .C(_3126__bF_buf6), .Y(_4656_) );
	AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_4645_), .B(_3126__bF_buf5), .C(_4656_), .Y(_4657_) );
	OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf0), .B(_4657_), .C(_4633_), .Y(csr_gpr_iu_rs1_27_) );
	NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__28_), .B(_3113__bF_buf15), .C(_3111__bF_buf15), .Y(_4658_) );
	MUX2X1 MUX2X1_84 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__28_), .B(csr_gpr_iu_gpr_29__28_), .S(biu_ins_15_bF_buf4), .Y(_4659_) );
	OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_4659_), .B(_3127__bF_buf1), .C(_4658_), .Y(_4660_) );
	NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf0), .B(_4660_), .Y(_4661_) );
	INVX1 INVX1_1017 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__28_), .Y(_4662_) );
	NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__28_), .B(_3095__bF_buf11), .Y(_4663_) );
	OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_3113__bF_buf14), .C(_4663_), .Y(_4664_) );
	INVX1 INVX1_1018 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__28_), .Y(_4665_) );
	INVX1 INVX1_1019 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__28_), .Y(_4666_) );
	OAI22X1 OAI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(_4666_), .B(_3110__bF_buf11), .C(_4665_), .D(_3111__bF_buf14), .Y(_4667_) );
	OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(_4664_), .C(_3117__bF_buf6), .Y(_4668_) );
	NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf4), .B(_4668_), .C(_4661_), .Y(_4669_) );
	OAI22X1 OAI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .B(_3110__bF_buf10), .C(_2853_), .D(_3111__bF_buf13), .Y(_4670_) );
	NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__28_), .B(_3095__bF_buf10), .Y(_4671_) );
	OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_3113__bF_buf13), .C(_4671_), .Y(_4672_) );
	OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .B(_4672_), .C(_3109__bF_buf10), .Y(_4673_) );
	INVX1 INVX1_1020 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__28_), .Y(_4674_) );
	OAI22X1 OAI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3110__bF_buf9), .C(_4674_), .D(_3111__bF_buf12), .Y(_4675_) );
	INVX1 INVX1_1021 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__28_), .Y(_4676_) );
	NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__28_), .B(_3095__bF_buf9), .Y(_4677_) );
	OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_3113__bF_buf12), .C(_4677_), .Y(_4678_) );
	OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_4675_), .B(_4678_), .C(_3117__bF_buf5), .Y(_4679_) );
	NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_4679_), .C(_3107__bF_buf1), .Y(_4680_) );
	NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4680_), .C(_4669_), .Y(_4681_) );
	INVX1 INVX1_1022 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__28_), .Y(_4682_) );
	INVX1 INVX1_1023 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__28_), .Y(_4683_) );
	OAI22X1 OAI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_3110__bF_buf8), .C(_4682_), .D(_3111__bF_buf11), .Y(_4684_) );
	INVX1 INVX1_1024 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__28_), .Y(_4685_) );
	NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__28_), .B(_3095__bF_buf8), .Y(_4686_) );
	OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_4685_), .B(_3113__bF_buf11), .C(_4686_), .Y(_4687_) );
	OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_4687_), .C(_3109__bF_buf9), .Y(_4688_) );
	INVX1 INVX1_1025 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__28_), .Y(_4689_) );
	NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__28_), .B(_3095__bF_buf7), .Y(_4690_) );
	OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_4689_), .B(_3113__bF_buf10), .C(_4690_), .Y(_4691_) );
	INVX1 INVX1_1026 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__28_), .Y(_4692_) );
	INVX1 INVX1_1027 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__28_), .Y(_4693_) );
	OAI22X1 OAI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_3110__bF_buf7), .C(_4692_), .D(_3111__bF_buf10), .Y(_4694_) );
	OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(_4691_), .C(_3117__bF_buf4), .Y(_4695_) );
	AOI22X1 AOI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4688_), .D(_4695_), .Y(_4696_) );
	INVX1 INVX1_1028 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__28_), .Y(_4697_) );
	INVX1 INVX1_1029 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__28_), .Y(_4698_) );
	OAI22X1 OAI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_3110__bF_buf6), .C(_4697_), .D(_3111__bF_buf9), .Y(_4699_) );
	INVX1 INVX1_1030 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__28_), .Y(_4700_) );
	NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__28_), .B(_3095__bF_buf6), .Y(_4701_) );
	OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(_3113__bF_buf9), .C(_4701_), .Y(_4702_) );
	OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_4699_), .B(_4702_), .C(_3109__bF_buf8), .Y(_4703_) );
	INVX1 INVX1_1031 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__28_), .Y(_4704_) );
	INVX1 INVX1_1032 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__28_), .Y(_4705_) );
	OAI22X1 OAI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4705_), .B(_3110__bF_buf5), .C(_4704_), .D(_3111__bF_buf8), .Y(_4706_) );
	INVX1 INVX1_1033 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__28_), .Y(_4707_) );
	NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__28_), .B(_3095__bF_buf5), .Y(_4708_) );
	OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_4707_), .B(_3113__bF_buf8), .C(_4708_), .Y(_4709_) );
	OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_4709_), .C(_3117__bF_buf3), .Y(_4710_) );
	AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_4703_), .B(_4710_), .C(_3107__bF_buf0), .Y(_4711_) );
	OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_4696_), .B(_4711_), .C(_3156__bF_buf1), .Y(_4712_) );
	AOI22X1 AOI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4681_), .D(_4712_), .Y(csr_gpr_iu_rs1_28_) );
	NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__29_), .B(_3113__bF_buf7), .C(_3111__bF_buf7), .Y(_4713_) );
	MUX2X1 MUX2X1_85 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__29_), .B(csr_gpr_iu_gpr_29__29_), .S(biu_ins_15_bF_buf3), .Y(_4714_) );
	OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .B(_3127__bF_buf0), .C(_4713_), .Y(_4715_) );
	NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3109__bF_buf7), .B(_4715_), .Y(_4716_) );
	INVX1 INVX1_1034 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__29_), .Y(_4717_) );
	INVX1 INVX1_1035 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__29_), .Y(_4718_) );
	OAI22X1 OAI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_3113__bF_buf6), .C(_4717_), .D(_3105__bF_buf7), .Y(_4719_) );
	INVX1 INVX1_1036 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__29_), .Y(_4720_) );
	INVX1 INVX1_1037 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__29_), .Y(_4721_) );
	OAI22X1 OAI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_3110__bF_buf4), .C(_4720_), .D(_3111__bF_buf6), .Y(_4722_) );
	OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4719_), .C(_3117__bF_buf2), .Y(_4723_) );
	NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3126__bF_buf3), .B(_4723_), .C(_4716_), .Y(_4724_) );
	OAI22X1 OAI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_3110__bF_buf3), .C(_2855_), .D(_3111__bF_buf5), .Y(_4725_) );
	NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__29_), .B(_3095__bF_buf4), .Y(_4726_) );
	OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_3113__bF_buf5), .C(_4726_), .Y(_4727_) );
	OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_4725_), .B(_4727_), .C(_3109__bF_buf6), .Y(_4728_) );
	INVX1 INVX1_1038 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__29_), .Y(_4729_) );
	OAI22X1 OAI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_3110__bF_buf2), .C(_4729_), .D(_3111__bF_buf4), .Y(_4730_) );
	INVX1 INVX1_1039 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__29_), .Y(_4731_) );
	INVX1 INVX1_1040 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__29_), .Y(_4732_) );
	OAI22X1 OAI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(_3113__bF_buf4), .C(_4731_), .D(_3105__bF_buf6), .Y(_4733_) );
	OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_4730_), .B(_4733_), .C(_3117__bF_buf1), .Y(_4734_) );
	NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_4734_), .B(_4728_), .C(_3107__bF_buf5), .Y(_4735_) );
	NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_4735_), .C(_4724_), .Y(_4736_) );
	INVX1 INVX1_1041 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__29_), .Y(_4737_) );
	INVX1 INVX1_1042 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__29_), .Y(_4738_) );
	OAI22X1 OAI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_3110__bF_buf1), .C(_4737_), .D(_3111__bF_buf3), .Y(_4739_) );
	INVX1 INVX1_1043 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__29_), .Y(_4740_) );
	INVX1 INVX1_1044 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__29_), .Y(_4741_) );
	OAI22X1 OAI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_3113__bF_buf3), .C(_4741_), .D(_3105__bF_buf5), .Y(_4742_) );
	OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_4739_), .B(_4742_), .C(_3109__bF_buf5), .Y(_4743_) );
	INVX1 INVX1_1045 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__29_), .Y(_4744_) );
	INVX1 INVX1_1046 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__29_), .Y(_4745_) );
	OAI22X1 OAI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_3110__bF_buf0), .C(_4744_), .D(_3113__bF_buf2), .Y(_4746_) );
	INVX1 INVX1_1047 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__29_), .Y(_4747_) );
	INVX1 INVX1_1048 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__29_), .Y(_4748_) );
	OAI22X1 OAI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(_3111__bF_buf2), .C(_4748_), .D(_3105__bF_buf4), .Y(_4749_) );
	OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_4749_), .C(_3117__bF_buf0), .Y(_4750_) );
	AOI22X1 AOI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3106_), .C(_4743_), .D(_4750_), .Y(_4751_) );
	INVX1 INVX1_1049 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__29_), .Y(_4752_) );
	INVX1 INVX1_1050 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__29_), .Y(_4753_) );
	OAI22X1 OAI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_3111__bF_buf1), .C(_4753_), .D(_3105__bF_buf3), .Y(_4754_) );
	INVX1 INVX1_1051 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__29_), .Y(_4755_) );
	INVX1 INVX1_1052 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__29_), .Y(_4756_) );
	OAI22X1 OAI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_3110__bF_buf13), .C(_4755_), .D(_3113__bF_buf1), .Y(_4757_) );
	OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_4757_), .B(_4754_), .C(_3109__bF_buf4), .Y(_4758_) );
	INVX1 INVX1_1053 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__29_), .Y(_4759_) );
	INVX1 INVX1_1054 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__29_), .Y(_4760_) );
	OAI22X1 OAI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(_3111__bF_buf0), .C(_4760_), .D(_3105__bF_buf2), .Y(_4761_) );
	INVX1 INVX1_1055 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__29_), .Y(_4762_) );
	INVX1 INVX1_1056 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__29_), .Y(_4763_) );
	OAI22X1 OAI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_3110__bF_buf12), .C(_4762_), .D(_3113__bF_buf0), .Y(_4764_) );
	OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(_4761_), .C(_3117__bF_buf9), .Y(_4765_) );
	AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_4765_), .B(_4758_), .C(_3107__bF_buf4), .Y(_4766_) );
	OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_4751_), .B(_4766_), .C(_3156__bF_buf0), .Y(_4767_) );
	AOI22X1 AOI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3097_), .C(_4736_), .D(_4767_), .Y(csr_gpr_iu_rs1_29_) );
	INVX1 INVX1_1057 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__30_), .Y(_4768_) );
	INVX1 INVX1_1058 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__30_), .Y(_4769_) );
	OAI22X1 OAI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4769_), .B(_3110__bF_buf11), .C(_4768_), .D(_3105__bF_buf1), .Y(_4770_) );
	INVX1 INVX1_1059 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__30_), .Y(_4771_) );
	INVX1 INVX1_1060 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__30_), .Y(_4772_) );
	OAI22X1 OAI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(_4771_), .B(_3111__bF_buf15), .C(_4772_), .D(_3113__bF_buf15), .Y(_4773_) );
	OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4773_), .C(_3109__bF_buf3), .Y(_4774_) );
	INVX1 INVX1_1061 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__30_), .Y(_4775_) );
	INVX1 INVX1_1062 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__30_), .Y(_4776_) );
	OAI22X1 OAI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(_4776_), .B(_3110__bF_buf10), .C(_4775_), .D(_3105__bF_buf0), .Y(_4777_) );
	INVX1 INVX1_1063 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__30_), .Y(_4778_) );
	INVX1 INVX1_1064 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__30_), .Y(_4779_) );
	OAI22X1 OAI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_3111__bF_buf14), .C(_4779_), .D(_3113__bF_buf14), .Y(_4780_) );
	OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_4777_), .B(_4780_), .C(_3117__bF_buf8), .Y(_4781_) );
	AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(_4774_), .C(_3107__bF_buf3), .Y(_4782_) );
	INVX1 INVX1_1065 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__30_), .Y(_4783_) );
	INVX1 INVX1_1066 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__30_), .Y(_4784_) );
	OAI22X1 OAI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(_4784_), .B(_3110__bF_buf9), .C(_4783_), .D(_3113__bF_buf13), .Y(_4785_) );
	INVX1 INVX1_1067 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__30_), .Y(_4786_) );
	NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__30_), .B(_3095__bF_buf3), .Y(_4787_) );
	OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(_3111__bF_buf13), .C(_4787_), .Y(_4788_) );
	OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_4788_), .C(_3109__bF_buf2), .Y(_4789_) );
	INVX1 INVX1_1068 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__30_), .Y(_4790_) );
	INVX1 INVX1_1069 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__30_), .Y(_4791_) );
	OAI22X1 OAI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(_4791_), .B(_3110__bF_buf8), .C(_4790_), .D(_3113__bF_buf12), .Y(_4792_) );
	INVX1 INVX1_1070 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__30_), .Y(_4793_) );
	NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__30_), .B(_3095__bF_buf2), .Y(_4794_) );
	OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(_3111__bF_buf12), .C(_4794_), .Y(_4795_) );
	OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_4795_), .C(_3117__bF_buf7), .Y(_4796_) );
	AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(_4796_), .C(_3126__bF_buf2), .Y(_4797_) );
	OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_4782_), .B(_4797_), .C(_3156__bF_buf4), .Y(_4798_) );
	INVX1 INVX1_1071 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__30_), .Y(_4799_) );
	INVX1 INVX1_1072 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__30_), .Y(_4800_) );
	OAI22X1 OAI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4799_), .B(_3111__bF_buf11), .C(_4800_), .D(_3113__bF_buf11), .Y(_4801_) );
	INVX1 INVX1_1073 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__30_), .Y(_4802_) );
	NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__30_), .B(biu_ins_15_bF_buf2), .Y(_4803_) );
	OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf1), .B(_4802_), .C(_4803_), .Y(_4804_) );
	AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf5), .B(_4804_), .C(_4801_), .Y(_4805_) );
	INVX1 INVX1_1074 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__30_), .Y(_4806_) );
	INVX1 INVX1_1075 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__30_), .Y(_4807_) );
	OAI22X1 OAI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(_3111__bF_buf10), .C(_4807_), .D(_3113__bF_buf10), .Y(_4808_) );
	AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__30_), .B(_3127__bF_buf4), .C(_4808_), .Y(_4809_) );
	MUX2X1 MUX2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_4805_), .S(_3109__bF_buf1), .Y(_4810_) );
	NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__30_), .B(_3095__bF_buf1), .Y(_4811_) );
	OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_3111__bF_buf9), .C(_4811_), .Y(_4812_) );
	OAI22X1 OAI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_3110__bF_buf7), .C(_2792_), .D(_3113__bF_buf9), .Y(_4813_) );
	OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4812_), .C(_3109__bF_buf0), .Y(_4814_) );
	INVX1 INVX1_1076 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__30_), .Y(_4815_) );
	INVX1 INVX1_1077 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__30_), .Y(_4816_) );
	OAI22X1 OAI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_3111__bF_buf8), .C(_4816_), .D(_3113__bF_buf8), .Y(_4817_) );
	INVX1 INVX1_1078 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__30_), .Y(_4818_) );
	OAI22X1 OAI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3110__bF_buf6), .C(_4818_), .D(_3105__bF_buf7), .Y(_4819_) );
	OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(_4817_), .C(_3117__bF_buf6), .Y(_4820_) );
	AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_4814_), .B(_4820_), .C(_3126__bF_buf1), .Y(_4821_) );
	AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_4810_), .B(_3126__bF_buf0), .C(_4821_), .Y(_4822_) );
	OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf3), .B(_4822_), .C(_4798_), .Y(csr_gpr_iu_rs1_30_) );
	INVX1 INVX1_1079 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__31_), .Y(_4823_) );
	INVX1 INVX1_1080 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_14__31_), .Y(_4824_) );
	OAI22X1 OAI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_3110__bF_buf5), .C(_4823_), .D(_3105__bF_buf6), .Y(_4825_) );
	INVX1 INVX1_1081 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_13__31_), .Y(_4826_) );
	INVX1 INVX1_1082 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_12__31_), .Y(_4827_) );
	OAI22X1 OAI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_3111__bF_buf7), .C(_4827_), .D(_3113__bF_buf7), .Y(_4828_) );
	OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_4825_), .B(_4828_), .C(_3109__bF_buf10), .Y(_4829_) );
	INVX1 INVX1_1083 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__31_), .Y(_4830_) );
	INVX1 INVX1_1084 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_10__31_), .Y(_4831_) );
	OAI22X1 OAI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(_4831_), .B(_3110__bF_buf4), .C(_4830_), .D(_3105__bF_buf5), .Y(_4832_) );
	INVX1 INVX1_1085 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_9__31_), .Y(_4833_) );
	INVX1 INVX1_1086 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_8__31_), .Y(_4834_) );
	OAI22X1 OAI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_3111__bF_buf6), .C(_4834_), .D(_3113__bF_buf6), .Y(_4835_) );
	OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_4835_), .C(_3117__bF_buf5), .Y(_4836_) );
	AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_4836_), .B(_4829_), .C(_3107__bF_buf2), .Y(_4837_) );
	INVX1 INVX1_1087 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_4__31_), .Y(_4838_) );
	INVX1 INVX1_1088 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__31_), .Y(_4839_) );
	OAI22X1 OAI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .B(_3113__bF_buf5), .C(_4839_), .D(_3105__bF_buf4), .Y(_4840_) );
	INVX1 INVX1_1089 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_5__31_), .Y(_4841_) );
	INVX1 INVX1_1090 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_6__31_), .Y(_4842_) );
	OAI22X1 OAI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_3110__bF_buf3), .C(_4841_), .D(_3111__bF_buf5), .Y(_4843_) );
	OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(_4840_), .C(_3109__bF_buf9), .Y(_4844_) );
	INVX1 INVX1_1091 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_0__31_), .Y(_4845_) );
	INVX1 INVX1_1092 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__31_), .Y(_4846_) );
	OAI22X1 OAI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(_4845_), .B(_3113__bF_buf4), .C(_4846_), .D(_3105__bF_buf3), .Y(_4847_) );
	INVX1 INVX1_1093 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_1__31_), .Y(_4848_) );
	INVX1 INVX1_1094 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_2__31_), .Y(_4849_) );
	OAI22X1 OAI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .B(_3110__bF_buf2), .C(_4848_), .D(_3111__bF_buf4), .Y(_4850_) );
	OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .B(_4847_), .C(_3117__bF_buf4), .Y(_4851_) );
	AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(_4844_), .C(_3126__bF_buf7), .Y(_4852_) );
	OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_4837_), .B(_4852_), .C(_3156__bF_buf3), .Y(_4853_) );
	INVX1 INVX1_1095 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_25__31_), .Y(_4854_) );
	INVX1 INVX1_1096 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_24__31_), .Y(_4855_) );
	OAI22X1 OAI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(_4854_), .B(_3111__bF_buf3), .C(_4855_), .D(_3113__bF_buf3), .Y(_4856_) );
	INVX1 INVX1_1097 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__31_), .Y(_4857_) );
	NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__31_), .B(biu_ins_15_bF_buf0), .Y(_4858_) );
	OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf6), .B(_4857_), .C(_4858_), .Y(_4859_) );
	AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3127__bF_buf3), .B(_4859_), .C(_4856_), .Y(_4860_) );
	INVX1 INVX1_1098 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__31_), .Y(_4861_) );
	INVX1 INVX1_1099 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__31_), .Y(_4862_) );
	OAI22X1 OAI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(_4861_), .B(_3111__bF_buf2), .C(_4862_), .D(_3113__bF_buf2), .Y(_4863_) );
	AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__31_), .B(_3127__bF_buf2), .C(_4863_), .Y(_4864_) );
	MUX2X1 MUX2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_4860_), .S(_3109__bF_buf8), .Y(_4865_) );
	NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__31_), .B(_3095__bF_buf0), .Y(_4866_) );
	OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_3111__bF_buf1), .C(_4866_), .Y(_4867_) );
	OAI22X1 OAI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_3110__bF_buf1), .C(_2794_), .D(_3113__bF_buf1), .Y(_4868_) );
	OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_4867_), .C(_3109__bF_buf7), .Y(_4869_) );
	INVX1 INVX1_1100 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_17__31_), .Y(_4870_) );
	INVX1 INVX1_1101 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_16__31_), .Y(_4871_) );
	OAI22X1 OAI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(_4870_), .B(_3111__bF_buf0), .C(_4871_), .D(_3113__bF_buf0), .Y(_4872_) );
	INVX1 INVX1_1102 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__31_), .Y(_4873_) );
	OAI22X1 OAI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .B(_3110__bF_buf0), .C(_4873_), .D(_3105__bF_buf2), .Y(_4874_) );
	OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_4874_), .B(_4872_), .C(_3117__bF_buf3), .Y(_4875_) );
	AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(_4875_), .C(_3126__bF_buf6), .Y(_4876_) );
	AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_3126__bF_buf5), .C(_4876_), .Y(_4877_) );
	OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_3100__bF_buf2), .B(_4877_), .C(_4853_), .Y(csr_gpr_iu_rs1_31_) );
	INVX8 INVX8_50 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_4878_) );
	INVX1 INVX1_1103 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf2), .Y(_4879_) );
	INVX1 INVX1_1104 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .Y(_4880_) );
	NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf5), .B(biu_ins_21_bF_buf2), .Y(_4881_) );
	NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_4879_), .B(_4880_), .C(_4881__bF_buf11), .Y(_4882_) );
	INVX8 INVX8_51 ( .gnd(gnd), .vdd(vdd), .A(_4882_), .Y(_4883_) );
	NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .Y(_4884_) );
	NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_4879_), .B(_4881__bF_buf10), .Y(_4885_) );
	OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .B(_4885_), .C(biu_ins_24_), .Y(_4886_) );
	NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf3), .B(_4884_), .Y(_4887_) );
	OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_4885_), .B(_4880_), .Y(_4888_) );
	INVX1 INVX1_1105 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf4), .Y(_4889_) );
	INVX1 INVX1_1106 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf1), .Y(_4890_) );
	NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4889_), .B(_4890_), .Y(_4891_) );
	OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf1), .B(_4891__bF_buf7), .C(_4880_), .Y(_4892_) );
	NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_4888_), .Y(_4893_) );
	OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(biu_ins_21_bF_buf0), .C(biu_ins_22_bF_buf0), .Y(_4894_) );
	NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4894_), .B(_4885_), .Y(_4895_) );
	NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf2), .B(biu_ins_21_bF_buf3), .Y(_4896_) );
	NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf2), .B(_4889_), .Y(_4897_) );
	OAI22X1 OAI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_4896__bF_buf13), .C(_2796_), .D(_4897__bF_buf15), .Y(_4898_) );
	NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf1), .B(_4890_), .Y(_4899_) );
	NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__0_), .B(_4881__bF_buf9), .Y(_4900_) );
	OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_2729_), .B(_4899__bF_buf15), .C(_4900_), .Y(_4901_) );
	OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_4901_), .C(_4895__bF_buf10), .Y(_4902_) );
	AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_4885_), .B(_4894_), .Y(_4903_) );
	OAI22X1 OAI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_4896__bF_buf12), .C(_3118_), .D(_4897__bF_buf14), .Y(_4904_) );
	NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__0_), .B(_4881__bF_buf8), .Y(_4905_) );
	OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_4899__bF_buf14), .C(_4905_), .Y(_4906_) );
	OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_4904_), .B(_4906_), .C(_4903__bF_buf9), .Y(_4907_) );
	NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_4902_), .B(_4907_), .C(_4893__bF_buf5), .Y(_4908_) );
	OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf3), .B(_4891__bF_buf6), .C(biu_ins_23_), .Y(_4909_) );
	NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_4882_), .B(_4909_), .Y(_4910_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf0), .B(biu_ins_21_bF_buf1), .Y(_4911_) );
	NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__0_), .B(_4899__bF_buf13), .C(_4897__bF_buf13), .Y(_4912_) );
	MUX2X1 MUX2X1_88 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__0_), .B(csr_gpr_iu_gpr_29__0_), .S(biu_ins_20_bF_buf6), .Y(_4913_) );
	OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_4913_), .B(_4911__bF_buf5), .C(_4912_), .Y(_4914_) );
	NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf9), .B(_4914_), .Y(_4915_) );
	NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__0_), .B(_4881__bF_buf7), .Y(_4916_) );
	OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_3132_), .B(_4899__bF_buf12), .C(_4916_), .Y(_4917_) );
	OAI22X1 OAI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_4896__bF_buf11), .C(_3135_), .D(_4897__bF_buf12), .Y(_4918_) );
	OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_4918_), .B(_4917_), .C(_4903__bF_buf8), .Y(_4919_) );
	NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_4919_), .C(_4915_), .Y(_4920_) );
	NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_4908_), .C(_4920_), .Y(_4921_) );
	OAI22X1 OAI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_4896__bF_buf10), .C(_3160_), .D(_4897__bF_buf11), .Y(_4922_) );
	NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__0_), .B(_4881__bF_buf6), .Y(_4923_) );
	OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .B(_4899__bF_buf11), .C(_4923_), .Y(_4924_) );
	OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_4922_), .B(_4924_), .C(_4895__bF_buf8), .Y(_4925_) );
	OAI22X1 OAI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(_3168_), .B(_4896__bF_buf9), .C(_3164_), .D(_4899__bF_buf10), .Y(_4926_) );
	NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__0_), .B(_4881__bF_buf5), .Y(_4927_) );
	OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_3167_), .B(_4897__bF_buf10), .C(_4927_), .Y(_4928_) );
	OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_4926_), .B(_4928_), .C(_4903__bF_buf7), .Y(_4929_) );
	AOI22X1 AOI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_4925_), .D(_4929_), .Y(_4930_) );
	INVX8 INVX8_52 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .Y(_4931_) );
	NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__0_), .B(_4881__bF_buf4), .Y(_4932_) );
	OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_4897__bF_buf9), .C(_4932_), .Y(_4933_) );
	OAI22X1 OAI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(_3142_), .B(_4896__bF_buf8), .C(_3141_), .D(_4899__bF_buf9), .Y(_4934_) );
	OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_4933_), .C(_4895__bF_buf7), .Y(_4935_) );
	NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__0_), .B(_4881__bF_buf3), .Y(_4936_) );
	OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_4897__bF_buf8), .C(_4936_), .Y(_4937_) );
	OAI22X1 OAI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_4896__bF_buf7), .C(_3151_), .D(_4899__bF_buf8), .Y(_4938_) );
	OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(_4937_), .C(_4903__bF_buf6), .Y(_4939_) );
	AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_4939_), .C(_4893__bF_buf4), .Y(_4940_) );
	OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4940_), .C(_4931__bF_buf4), .Y(_4941_) );
	AOI22X1 AOI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_4921_), .D(_4941_), .Y(csr_gpr_iu_rs2_0_) );
	NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__1_), .B(_4899__bF_buf7), .C(_4897__bF_buf7), .Y(_4942_) );
	MUX2X1 MUX2X1_89 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__1_), .B(csr_gpr_iu_gpr_29__1_), .S(biu_ins_20_bF_buf5), .Y(_4943_) );
	OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4911__bF_buf4), .C(_4942_), .Y(_4944_) );
	NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf6), .B(_4944_), .Y(_4945_) );
	NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__1_), .B(_4881__bF_buf2), .Y(_4946_) );
	OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_4899__bF_buf6), .C(_4946_), .Y(_4947_) );
	OAI22X1 OAI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(_3181_), .B(_4896__bF_buf6), .C(_3180_), .D(_4897__bF_buf6), .Y(_4948_) );
	OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_4948_), .B(_4947_), .C(_4903__bF_buf5), .Y(_4949_) );
	NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf6), .B(_4949_), .C(_4945_), .Y(_4950_) );
	OAI22X1 OAI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_4896__bF_buf5), .C(_2799_), .D(_4897__bF_buf5), .Y(_4951_) );
	NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__1_), .B(_4881__bF_buf1), .Y(_4952_) );
	OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_4899__bF_buf5), .C(_4952_), .Y(_4953_) );
	OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_4951_), .B(_4953_), .C(_4895__bF_buf5), .Y(_4954_) );
	OAI22X1 OAI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_4896__bF_buf4), .C(_3189_), .D(_4897__bF_buf4), .Y(_4955_) );
	NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__1_), .B(_4881__bF_buf0), .Y(_4956_) );
	OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .B(_4899__bF_buf4), .C(_4956_), .Y(_4957_) );
	OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4957_), .C(_4903__bF_buf4), .Y(_4958_) );
	NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_4954_), .B(_4958_), .C(_4893__bF_buf3), .Y(_4959_) );
	NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_4959_), .C(_4950_), .Y(_4960_) );
	NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__1_), .B(_4881__bF_buf11), .Y(_4961_) );
	OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(_4897__bF_buf3), .C(_4961_), .Y(_4962_) );
	OAI22X1 OAI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_4896__bF_buf3), .C(_3200_), .D(_4899__bF_buf3), .Y(_4963_) );
	OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4962_), .C(_4895__bF_buf4), .Y(_4964_) );
	OAI22X1 OAI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(_3205_), .B(_4896__bF_buf2), .C(_3204_), .D(_4899__bF_buf2), .Y(_4965_) );
	NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__1_), .B(_4881__bF_buf10), .Y(_4966_) );
	OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .B(_4897__bF_buf2), .C(_4966_), .Y(_4967_) );
	OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_4965_), .B(_4967_), .C(_4903__bF_buf3), .Y(_4968_) );
	AOI22X1 AOI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_4964_), .D(_4968_), .Y(_4969_) );
	OAI22X1 OAI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_4896__bF_buf1), .C(_3212_), .D(_4897__bF_buf1), .Y(_4970_) );
	NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__1_), .B(_4881__bF_buf9), .Y(_4971_) );
	OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_4899__bF_buf1), .C(_4971_), .Y(_4972_) );
	OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_4970_), .B(_4972_), .C(_4895__bF_buf3), .Y(_4973_) );
	OAI22X1 OAI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(_3220_), .B(_4896__bF_buf0), .C(_3219_), .D(_4897__bF_buf0), .Y(_4974_) );
	NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__1_), .B(_4881__bF_buf8), .Y(_4975_) );
	OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_4899__bF_buf0), .C(_4975_), .Y(_4976_) );
	OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .B(_4976_), .C(_4903__bF_buf2), .Y(_4977_) );
	AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .B(_4977_), .C(_4893__bF_buf2), .Y(_4978_) );
	OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_4969_), .B(_4978_), .C(_4931__bF_buf3), .Y(_4979_) );
	AOI22X1 AOI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_4960_), .D(_4979_), .Y(csr_gpr_iu_rs2_1_) );
	OAI22X1 OAI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(_3229_), .B(_4896__bF_buf13), .C(_3228_), .D(_4891__bF_buf5), .Y(_4980_) );
	OAI22X1 OAI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_4897__bF_buf15), .C(_3232_), .D(_4899__bF_buf15), .Y(_4981_) );
	OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .B(_4981_), .C(_4895__bF_buf2), .Y(_4982_) );
	OAI22X1 OAI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_4896__bF_buf12), .C(_3235_), .D(_4891__bF_buf4), .Y(_4983_) );
	OAI22X1 OAI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_4897__bF_buf14), .C(_3239_), .D(_4899__bF_buf14), .Y(_4984_) );
	OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(_4984_), .C(_4903__bF_buf1), .Y(_4985_) );
	AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_4985_), .B(_4982_), .C(_4893__bF_buf1), .Y(_4986_) );
	OAI22X1 OAI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_4896__bF_buf11), .C(_3244_), .D(_4899__bF_buf13), .Y(_4987_) );
	NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__2_), .B(_4881__bF_buf7), .Y(_4988_) );
	OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_4897__bF_buf13), .C(_4988_), .Y(_4989_) );
	OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_4989_), .C(_4895__bF_buf1), .Y(_4990_) );
	OAI22X1 OAI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_4896__bF_buf10), .C(_3251_), .D(_4899__bF_buf12), .Y(_4991_) );
	NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__2_), .B(_4881__bF_buf6), .Y(_4992_) );
	OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_4897__bF_buf12), .C(_4992_), .Y(_4993_) );
	OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_4991_), .B(_4993_), .C(_4903__bF_buf0), .Y(_4994_) );
	AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .B(_4994_), .C(_4910__bF_buf5), .Y(_4995_) );
	OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_4986_), .B(_4995_), .C(_4931__bF_buf2), .Y(_4996_) );
	OAI22X1 OAI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_4897__bF_buf11), .C(_3260_), .D(_4899__bF_buf11), .Y(_4997_) );
	NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__2_), .B(biu_ins_20_bF_buf4), .Y(_4998_) );
	OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(_3262_), .C(_4998_), .Y(_4999_) );
	AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf3), .B(_4999_), .C(_4997_), .Y(_5000_) );
	OAI22X1 OAI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .B(_4897__bF_buf10), .C(_3267_), .D(_4899__bF_buf10), .Y(_5001_) );
	AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__2_), .B(_4911__bF_buf2), .C(_5001_), .Y(_5002_) );
	MUX2X1 MUX2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_5002_), .B(_5000_), .S(_4895__bF_buf0), .Y(_5003_) );
	OAI22X1 OAI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_4896__bF_buf9), .C(_2801_), .D(_4897__bF_buf9), .Y(_5004_) );
	NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__2_), .B(_4881__bF_buf5), .Y(_5005_) );
	OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(_4899__bF_buf9), .C(_5005_), .Y(_5006_) );
	OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_5006_), .C(_4895__bF_buf10), .Y(_5007_) );
	OAI22X1 OAI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_4897__bF_buf8), .C(_3276_), .D(_4899__bF_buf8), .Y(_5008_) );
	OAI22X1 OAI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_4896__bF_buf8), .C(_3278_), .D(_4891__bF_buf3), .Y(_5009_) );
	OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_5009_), .B(_5008_), .C(_4903__bF_buf9), .Y(_5010_) );
	AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_5007_), .B(_5010_), .C(_4910__bF_buf4), .Y(_5011_) );
	AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_5003_), .B(_4910__bF_buf3), .C(_5011_), .Y(_5012_) );
	OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf2), .B(_5012_), .C(_4996_), .Y(csr_gpr_iu_rs2_2_) );
	OAI22X1 OAI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_4896__bF_buf7), .C(_3283_), .D(_4891__bF_buf2), .Y(_5013_) );
	OAI22X1 OAI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_4897__bF_buf7), .C(_3287_), .D(_4899__bF_buf7), .Y(_5014_) );
	OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_5013_), .B(_5014_), .C(_4895__bF_buf9), .Y(_5015_) );
	OAI22X1 OAI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(_3291_), .B(_4896__bF_buf6), .C(_3290_), .D(_4891__bF_buf1), .Y(_5016_) );
	OAI22X1 OAI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_4897__bF_buf6), .C(_3294_), .D(_4899__bF_buf6), .Y(_5017_) );
	OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(_5017_), .C(_4903__bF_buf8), .Y(_5018_) );
	AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_5018_), .B(_5015_), .C(_4893__bF_buf0), .Y(_5019_) );
	OAI22X1 OAI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(_3301_), .B(_4897__bF_buf5), .C(_3298_), .D(_4899__bF_buf5), .Y(_5020_) );
	OAI22X1 OAI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_4896__bF_buf5), .C(_3302_), .D(_4891__bF_buf0), .Y(_5021_) );
	OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_5020_), .C(_4895__bF_buf8), .Y(_5022_) );
	OAI22X1 OAI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_4897__bF_buf4), .C(_3305_), .D(_4899__bF_buf4), .Y(_5023_) );
	OAI22X1 OAI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_4896__bF_buf4), .C(_3309_), .D(_4891__bF_buf7), .Y(_5024_) );
	OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_5024_), .B(_5023_), .C(_4903__bF_buf7), .Y(_5025_) );
	AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5022_), .C(_4910__bF_buf2), .Y(_5026_) );
	OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(_5026_), .C(_4931__bF_buf1), .Y(_5027_) );
	OAI22X1 OAI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_4897__bF_buf3), .C(_3315_), .D(_4899__bF_buf3), .Y(_5028_) );
	NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__3_), .B(biu_ins_20_bF_buf2), .Y(_5029_) );
	OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf1), .B(_3317_), .C(_5029_), .Y(_5030_) );
	AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf1), .B(_5030_), .C(_5028_), .Y(_5031_) );
	OAI22X1 OAI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(_4897__bF_buf2), .C(_3322_), .D(_4899__bF_buf2), .Y(_5032_) );
	AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__3_), .B(_4911__bF_buf0), .C(_5032_), .Y(_5033_) );
	MUX2X1 MUX2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_5033_), .B(_5031_), .S(_4895__bF_buf7), .Y(_5034_) );
	NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__3_), .B(_4881__bF_buf4), .Y(_5035_) );
	OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_4897__bF_buf1), .C(_5035_), .Y(_5036_) );
	OAI22X1 OAI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(_4896__bF_buf3), .C(_2738_), .D(_4899__bF_buf1), .Y(_5037_) );
	OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5036_), .C(_4895__bF_buf6), .Y(_5038_) );
	OAI22X1 OAI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_4897__bF_buf0), .C(_3331_), .D(_4899__bF_buf0), .Y(_5039_) );
	OAI22X1 OAI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(_4896__bF_buf2), .C(_3333_), .D(_4891__bF_buf6), .Y(_5040_) );
	OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_5039_), .C(_4903__bF_buf6), .Y(_5041_) );
	AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(_5041_), .C(_4910__bF_buf1), .Y(_5042_) );
	AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_5034_), .B(_4910__bF_buf0), .C(_5042_), .Y(_5043_) );
	OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf1), .B(_5043_), .C(_5027_), .Y(csr_gpr_iu_rs2_3_) );
	NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__4_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5044_) );
	MUX2X1 MUX2X1_92 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__4_), .B(csr_gpr_iu_gpr_29__4_), .S(biu_ins_20_bF_buf0), .Y(_5045_) );
	OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_5045_), .B(_4911__bF_buf5), .C(_5044_), .Y(_5046_) );
	NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf5), .B(_5046_), .Y(_5047_) );
	NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__4_), .B(_4881__bF_buf3), .Y(_5048_) );
	OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .B(_4899__bF_buf14), .C(_5048_), .Y(_5049_) );
	OAI22X1 OAI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_4896__bF_buf1), .C(_3345_), .D(_4897__bF_buf14), .Y(_5050_) );
	OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_5050_), .B(_5049_), .C(_4903__bF_buf5), .Y(_5051_) );
	NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_5051_), .C(_5047_), .Y(_5052_) );
	NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__4_), .B(_4881__bF_buf2), .Y(_5053_) );
	OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_4897__bF_buf13), .C(_5053_), .Y(_5054_) );
	OAI22X1 OAI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_4896__bF_buf0), .C(_2740_), .D(_4899__bF_buf13), .Y(_5055_) );
	OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_5054_), .C(_4895__bF_buf4), .Y(_5056_) );
	NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__4_), .B(_4881__bF_buf1), .Y(_5057_) );
	OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(_4897__bF_buf12), .C(_5057_), .Y(_5058_) );
	OAI22X1 OAI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_4896__bF_buf13), .C(_3357_), .D(_4899__bF_buf12), .Y(_5059_) );
	OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(_5058_), .C(_4903__bF_buf4), .Y(_5060_) );
	NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_5056_), .B(_5060_), .C(_4893__bF_buf5), .Y(_5061_) );
	NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5061_), .C(_5052_), .Y(_5062_) );
	NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__4_), .B(_4881__bF_buf0), .Y(_5063_) );
	OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_4899__bF_buf11), .C(_5063_), .Y(_5064_) );
	OAI22X1 OAI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_4896__bF_buf12), .C(_3362_), .D(_4897__bF_buf11), .Y(_5065_) );
	OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_5065_), .B(_5064_), .C(_4895__bF_buf3), .Y(_5066_) );
	OAI22X1 OAI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_4896__bF_buf11), .C(_3372_), .D(_4897__bF_buf10), .Y(_5067_) );
	NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__4_), .B(_4881__bF_buf11), .Y(_5068_) );
	OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_4899__bF_buf10), .C(_5068_), .Y(_5069_) );
	OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_5069_), .C(_4903__bF_buf3), .Y(_5070_) );
	AOI22X1 AOI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5066_), .D(_5070_), .Y(_5071_) );
	OAI22X1 OAI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_4896__bF_buf10), .C(_3377_), .D(_4897__bF_buf9), .Y(_5072_) );
	NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__4_), .B(_4881__bF_buf10), .Y(_5073_) );
	OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_3380_), .B(_4899__bF_buf9), .C(_5073_), .Y(_5074_) );
	OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_5072_), .B(_5074_), .C(_4895__bF_buf2), .Y(_5075_) );
	OAI22X1 OAI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_4896__bF_buf9), .C(_3384_), .D(_4897__bF_buf8), .Y(_5076_) );
	NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__4_), .B(_4881__bF_buf9), .Y(_5077_) );
	OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(_4899__bF_buf8), .C(_5077_), .Y(_5078_) );
	OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .B(_5078_), .C(_4903__bF_buf2), .Y(_5079_) );
	AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_5079_), .C(_4893__bF_buf4), .Y(_5080_) );
	OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_5071_), .B(_5080_), .C(_4931__bF_buf0), .Y(_5081_) );
	AOI22X1 AOI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5062_), .D(_5081_), .Y(csr_gpr_iu_rs2_4_) );
	OAI22X1 OAI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3394_), .B(_4896__bF_buf8), .C(_3393_), .D(_4891__bF_buf5), .Y(_5082_) );
	OAI22X1 OAI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_4897__bF_buf7), .C(_3397_), .D(_4899__bF_buf7), .Y(_5083_) );
	OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5083_), .C(_4895__bF_buf1), .Y(_5084_) );
	OAI22X1 OAI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(_3401_), .B(_4896__bF_buf7), .C(_3400_), .D(_4891__bF_buf4), .Y(_5085_) );
	OAI22X1 OAI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_4897__bF_buf6), .C(_3404_), .D(_4899__bF_buf6), .Y(_5086_) );
	OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .B(_5086_), .C(_4903__bF_buf1), .Y(_5087_) );
	AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5084_), .C(_4893__bF_buf3), .Y(_5088_) );
	NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__5_), .B(_4881__bF_buf8), .Y(_5089_) );
	OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_4899__bF_buf5), .C(_5089_), .Y(_5090_) );
	OAI22X1 OAI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_4896__bF_buf6), .C(_3411_), .D(_4897__bF_buf5), .Y(_5091_) );
	OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .B(_5090_), .C(_4895__bF_buf0), .Y(_5092_) );
	NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__5_), .B(_4881__bF_buf7), .Y(_5093_) );
	OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_3415_), .B(_4899__bF_buf4), .C(_5093_), .Y(_5094_) );
	OAI22X1 OAI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_4896__bF_buf5), .C(_3418_), .D(_4897__bF_buf4), .Y(_5095_) );
	OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5094_), .C(_4903__bF_buf0), .Y(_5096_) );
	AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .B(_5096_), .C(_4910__bF_buf6), .Y(_5097_) );
	OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5097_), .C(_4931__bF_buf4), .Y(_5098_) );
	OAI22X1 OAI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(_3424_), .B(_4897__bF_buf3), .C(_3425_), .D(_4899__bF_buf3), .Y(_5099_) );
	NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__5_), .B(biu_ins_20_bF_buf6), .Y(_5100_) );
	OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf5), .B(_3427_), .C(_5100_), .Y(_5101_) );
	AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf4), .B(_5101_), .C(_5099_), .Y(_5102_) );
	OAI22X1 OAI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .B(_4897__bF_buf2), .C(_3432_), .D(_4899__bF_buf2), .Y(_5103_) );
	AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__5_), .B(_4911__bF_buf3), .C(_5103_), .Y(_5104_) );
	MUX2X1 MUX2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .B(_5102_), .S(_4895__bF_buf10), .Y(_5105_) );
	NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__5_), .B(_4881__bF_buf6), .Y(_5106_) );
	OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .B(_4897__bF_buf1), .C(_5106_), .Y(_5107_) );
	OAI22X1 OAI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_4896__bF_buf4), .C(_2742_), .D(_4899__bF_buf1), .Y(_5108_) );
	OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .B(_5107_), .C(_4895__bF_buf9), .Y(_5109_) );
	OAI22X1 OAI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_4897__bF_buf0), .C(_3441_), .D(_4899__bF_buf0), .Y(_5110_) );
	OAI22X1 OAI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_4896__bF_buf3), .C(_3443_), .D(_4891__bF_buf3), .Y(_5111_) );
	OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .B(_5110_), .C(_4903__bF_buf9), .Y(_5112_) );
	AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .B(_5112_), .C(_4910__bF_buf5), .Y(_5113_) );
	AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_4910__bF_buf4), .C(_5113_), .Y(_5114_) );
	OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf0), .B(_5114_), .C(_5098_), .Y(csr_gpr_iu_rs2_5_) );
	OAI22X1 OAI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_4896__bF_buf2), .C(_3448_), .D(_4891__bF_buf2), .Y(_5115_) );
	OAI22X1 OAI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_4897__bF_buf15), .C(_3452_), .D(_4899__bF_buf15), .Y(_5116_) );
	OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .B(_5116_), .C(_4895__bF_buf8), .Y(_5117_) );
	OAI22X1 OAI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(_3456_), .B(_4896__bF_buf1), .C(_3455_), .D(_4891__bF_buf1), .Y(_5118_) );
	OAI22X1 OAI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_4897__bF_buf14), .C(_3459_), .D(_4899__bF_buf14), .Y(_5119_) );
	OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .B(_5119_), .C(_4903__bF_buf8), .Y(_5120_) );
	AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .B(_5117_), .C(_4893__bF_buf2), .Y(_5121_) );
	OAI22X1 OAI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_4896__bF_buf0), .C(_3463_), .D(_4899__bF_buf13), .Y(_5122_) );
	NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__6_), .B(_4881__bF_buf5), .Y(_5123_) );
	OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_3466_), .B(_4897__bF_buf13), .C(_5123_), .Y(_5124_) );
	OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .B(_5124_), .C(_4895__bF_buf7), .Y(_5125_) );
	OAI22X1 OAI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(_4896__bF_buf13), .C(_3470_), .D(_4899__bF_buf12), .Y(_5126_) );
	NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__6_), .B(_4881__bF_buf4), .Y(_5127_) );
	OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_4897__bF_buf12), .C(_5127_), .Y(_5128_) );
	OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5128_), .C(_4903__bF_buf7), .Y(_5129_) );
	AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .B(_5129_), .C(_4910__bF_buf3), .Y(_5130_) );
	OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .B(_5130_), .C(_4931__bF_buf3), .Y(_5131_) );
	OAI22X1 OAI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_4897__bF_buf11), .C(_3480_), .D(_4899__bF_buf11), .Y(_5132_) );
	NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__6_), .B(biu_ins_20_bF_buf4), .Y(_5133_) );
	OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(_3482_), .C(_5133_), .Y(_5134_) );
	AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf2), .B(_5134_), .C(_5132_), .Y(_5135_) );
	OAI22X1 OAI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_4897__bF_buf10), .C(_3487_), .D(_4899__bF_buf10), .Y(_5136_) );
	AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__6_), .B(_4911__bF_buf1), .C(_5136_), .Y(_5137_) );
	MUX2X1 MUX2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_5137_), .B(_5135_), .S(_4895__bF_buf6), .Y(_5138_) );
	NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__6_), .B(_4881__bF_buf3), .Y(_5139_) );
	OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_2809_), .B(_4897__bF_buf9), .C(_5139_), .Y(_5140_) );
	OAI22X1 OAI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .B(_4896__bF_buf12), .C(_2744_), .D(_4899__bF_buf9), .Y(_5141_) );
	OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_5141_), .B(_5140_), .C(_4895__bF_buf5), .Y(_5142_) );
	OAI22X1 OAI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_4897__bF_buf8), .C(_3496_), .D(_4899__bF_buf8), .Y(_5143_) );
	OAI22X1 OAI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(_4896__bF_buf11), .C(_3498_), .D(_4891__bF_buf0), .Y(_5144_) );
	OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_5144_), .B(_5143_), .C(_4903__bF_buf6), .Y(_5145_) );
	AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_5145_), .C(_4910__bF_buf2), .Y(_5146_) );
	AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_5138_), .B(_4910__bF_buf1), .C(_5146_), .Y(_5147_) );
	OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf3), .B(_5147_), .C(_5131_), .Y(csr_gpr_iu_rs2_6_) );
	OAI22X1 OAI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_4896__bF_buf10), .C(_3543_), .D(_4891__bF_buf7), .Y(_5148_) );
	OAI22X1 OAI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_4897__bF_buf7), .C(_3545_), .D(_4899__bF_buf7), .Y(_5149_) );
	OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_5149_), .C(_4895__bF_buf4), .Y(_5150_) );
	OAI22X1 OAI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_4896__bF_buf9), .C(_3550_), .D(_4891__bF_buf6), .Y(_5151_) );
	OAI22X1 OAI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_4897__bF_buf6), .C(_3552_), .D(_4899__bF_buf6), .Y(_5152_) );
	OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_5151_), .B(_5152_), .C(_4903__bF_buf5), .Y(_5153_) );
	AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_5153_), .B(_5150_), .C(_4893__bF_buf1), .Y(_5154_) );
	OAI22X1 OAI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_4897__bF_buf5), .C(_3530_), .D(_4899__bF_buf5), .Y(_5155_) );
	OAI22X1 OAI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_4896__bF_buf8), .C(_3528_), .D(_4891__bF_buf5), .Y(_5156_) );
	OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_5156_), .B(_5155_), .C(_4895__bF_buf3), .Y(_5157_) );
	OAI22X1 OAI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(_4897__bF_buf4), .C(_3534_), .D(_4899__bF_buf4), .Y(_5158_) );
	OAI22X1 OAI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .B(_4896__bF_buf7), .C(_3535_), .D(_4891__bF_buf4), .Y(_5159_) );
	OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_5159_), .B(_5158_), .C(_4903__bF_buf4), .Y(_5160_) );
	AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5157_), .C(_4910__bF_buf0), .Y(_5161_) );
	OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5161_), .C(_4931__bF_buf2), .Y(_5162_) );
	INVX1 INVX1_1107 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__7_), .Y(_5163_) );
	INVX1 INVX1_1108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__7_), .Y(_5164_) );
	OAI22X1 OAI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_4897__bF_buf3), .C(_5164_), .D(_4899__bF_buf3), .Y(_5165_) );
	AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__7_), .B(_4911__bF_buf0), .C(_5165_), .Y(_5166_) );
	OAI22X1 OAI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_4899__bF_buf2), .C(_3507_), .D(_4891__bF_buf3), .Y(_5167_) );
	OAI22X1 OAI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_4896__bF_buf6), .C(_3510_), .D(_4897__bF_buf2), .Y(_5168_) );
	OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5168_), .C(_4903__bF_buf3), .Y(_5169_) );
	OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_4903__bF_buf2), .B(_5166_), .C(_5169_), .Y(_5170_) );
	NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__7_), .B(_4881__bF_buf2), .Y(_5171_) );
	OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_2811_), .B(_4897__bF_buf1), .C(_5171_), .Y(_5172_) );
	OAI22X1 OAI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_4896__bF_buf5), .C(_2746_), .D(_4899__bF_buf1), .Y(_5173_) );
	OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5172_), .C(_4895__bF_buf2), .Y(_5174_) );
	OAI22X1 OAI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_4897__bF_buf0), .C(_3522_), .D(_4899__bF_buf0), .Y(_5175_) );
	OAI22X1 OAI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_4896__bF_buf4), .C(_3519_), .D(_4891__bF_buf2), .Y(_5176_) );
	OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_5176_), .B(_5175_), .C(_4903__bF_buf1), .Y(_5177_) );
	AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_5177_), .C(_4910__bF_buf7), .Y(_5178_) );
	AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_5170_), .B(_4910__bF_buf6), .C(_5178_), .Y(_5179_) );
	OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf2), .B(_5179_), .C(_5162_), .Y(csr_gpr_iu_rs2_7_) );
	NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__8_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5180_) );
	MUX2X1 MUX2X1_95 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__8_), .B(csr_gpr_iu_gpr_29__8_), .S(biu_ins_20_bF_buf2), .Y(_5181_) );
	OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_5181_), .B(_4911__bF_buf5), .C(_5180_), .Y(_5182_) );
	NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf1), .B(_5182_), .Y(_5183_) );
	NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__8_), .B(_4881__bF_buf1), .Y(_5184_) );
	OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_4899__bF_buf14), .C(_5184_), .Y(_5185_) );
	OAI22X1 OAI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3566_), .B(_4896__bF_buf3), .C(_3565_), .D(_4897__bF_buf14), .Y(_5186_) );
	OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_5185_), .C(_4903__bF_buf0), .Y(_5187_) );
	NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf5), .B(_5187_), .C(_5183_), .Y(_5188_) );
	OAI22X1 OAI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_4896__bF_buf2), .C(_2813_), .D(_4897__bF_buf13), .Y(_5189_) );
	NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__8_), .B(_4881__bF_buf0), .Y(_5190_) );
	OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_4899__bF_buf13), .C(_5190_), .Y(_5191_) );
	OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_5189_), .B(_5191_), .C(_4895__bF_buf0), .Y(_5192_) );
	OAI22X1 OAI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3011_), .B(_4896__bF_buf1), .C(_3574_), .D(_4897__bF_buf12), .Y(_5193_) );
	NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__8_), .B(_4881__bF_buf11), .Y(_5194_) );
	OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .B(_4899__bF_buf12), .C(_5194_), .Y(_5195_) );
	OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_5193_), .B(_5195_), .C(_4903__bF_buf9), .Y(_5196_) );
	NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_5196_), .C(_4893__bF_buf0), .Y(_5197_) );
	NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5197_), .C(_5188_), .Y(_5198_) );
	OAI22X1 OAI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_4896__bF_buf0), .C(_3582_), .D(_4897__bF_buf11), .Y(_5199_) );
	NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__8_), .B(_4881__bF_buf10), .Y(_5200_) );
	OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_3585_), .B(_4899__bF_buf11), .C(_5200_), .Y(_5201_) );
	OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_5199_), .B(_5201_), .C(_4895__bF_buf10), .Y(_5202_) );
	OAI22X1 OAI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(_4896__bF_buf13), .C(_3589_), .D(_4899__bF_buf10), .Y(_5203_) );
	NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__8_), .B(_4881__bF_buf9), .Y(_5204_) );
	OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_3592_), .B(_4897__bF_buf10), .C(_5204_), .Y(_5205_) );
	OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_5203_), .B(_5205_), .C(_4903__bF_buf8), .Y(_5206_) );
	AOI22X1 AOI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5202_), .D(_5206_), .Y(_5207_) );
	OAI22X1 OAI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_4896__bF_buf12), .C(_3597_), .D(_4897__bF_buf9), .Y(_5208_) );
	NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__8_), .B(_4881__bF_buf8), .Y(_5209_) );
	OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_4899__bF_buf9), .C(_5209_), .Y(_5210_) );
	OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_5208_), .B(_5210_), .C(_4895__bF_buf9), .Y(_5211_) );
	OAI22X1 OAI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_4896__bF_buf11), .C(_3604_), .D(_4897__bF_buf8), .Y(_5212_) );
	NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__8_), .B(_4881__bF_buf7), .Y(_5213_) );
	OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .B(_4899__bF_buf8), .C(_5213_), .Y(_5214_) );
	OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_5212_), .B(_5214_), .C(_4903__bF_buf7), .Y(_5215_) );
	AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5215_), .C(_4893__bF_buf5), .Y(_5216_) );
	OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_5207_), .B(_5216_), .C(_4931__bF_buf1), .Y(_5217_) );
	AOI22X1 AOI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5198_), .D(_5217_), .Y(csr_gpr_iu_rs2_8_) );
	NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__9_), .B(_4899__bF_buf7), .C(_4897__bF_buf7), .Y(_5218_) );
	MUX2X1 MUX2X1_96 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__9_), .B(csr_gpr_iu_gpr_29__9_), .S(biu_ins_20_bF_buf1), .Y(_5219_) );
	OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .B(_4911__bF_buf4), .C(_5218_), .Y(_5220_) );
	NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf8), .B(_5220_), .Y(_5221_) );
	NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__9_), .B(_4881__bF_buf6), .Y(_5222_) );
	OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_4899__bF_buf6), .C(_5222_), .Y(_5223_) );
	OAI22X1 OAI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_4896__bF_buf10), .C(_3620_), .D(_4897__bF_buf6), .Y(_5224_) );
	OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_5224_), .B(_5223_), .C(_4903__bF_buf6), .Y(_5225_) );
	NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf4), .B(_5225_), .C(_5221_), .Y(_5226_) );
	OAI22X1 OAI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_4896__bF_buf9), .C(_2815_), .D(_4897__bF_buf5), .Y(_5227_) );
	NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__9_), .B(_4881__bF_buf5), .Y(_5228_) );
	OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_4899__bF_buf5), .C(_5228_), .Y(_5229_) );
	OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_5227_), .B(_5229_), .C(_4895__bF_buf7), .Y(_5230_) );
	OAI22X1 OAI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_4896__bF_buf8), .C(_3629_), .D(_4897__bF_buf4), .Y(_5231_) );
	NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__9_), .B(_4881__bF_buf4), .Y(_5232_) );
	OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_4899__bF_buf4), .C(_5232_), .Y(_5233_) );
	OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_5231_), .B(_5233_), .C(_4903__bF_buf5), .Y(_5234_) );
	NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(_5234_), .C(_4893__bF_buf4), .Y(_5235_) );
	NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5235_), .C(_5226_), .Y(_5236_) );
	NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__9_), .B(_4881__bF_buf3), .Y(_5237_) );
	OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_4897__bF_buf3), .C(_5237_), .Y(_5238_) );
	OAI22X1 OAI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_4896__bF_buf7), .C(_3640_), .D(_4899__bF_buf3), .Y(_5239_) );
	OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_5239_), .B(_5238_), .C(_4895__bF_buf6), .Y(_5240_) );
	OAI22X1 OAI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_4896__bF_buf6), .C(_3644_), .D(_4899__bF_buf2), .Y(_5241_) );
	NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__9_), .B(_4881__bF_buf2), .Y(_5242_) );
	OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_4897__bF_buf2), .C(_5242_), .Y(_5243_) );
	OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_5241_), .B(_5243_), .C(_4903__bF_buf4), .Y(_5244_) );
	AOI22X1 AOI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5240_), .D(_5244_), .Y(_5245_) );
	OAI22X1 OAI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(_3653_), .B(_4896__bF_buf5), .C(_3652_), .D(_4897__bF_buf1), .Y(_5246_) );
	NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__9_), .B(_4881__bF_buf1), .Y(_5247_) );
	OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(_4899__bF_buf1), .C(_5247_), .Y(_5248_) );
	OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_5246_), .B(_5248_), .C(_4895__bF_buf5), .Y(_5249_) );
	OAI22X1 OAI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_4896__bF_buf4), .C(_3659_), .D(_4897__bF_buf0), .Y(_5250_) );
	NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__9_), .B(_4881__bF_buf0), .Y(_5251_) );
	OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_4899__bF_buf0), .C(_5251_), .Y(_5252_) );
	OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_5250_), .B(_5252_), .C(_4903__bF_buf3), .Y(_5253_) );
	AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(_5253_), .C(_4893__bF_buf3), .Y(_5254_) );
	OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_5245_), .B(_5254_), .C(_4931__bF_buf0), .Y(_5255_) );
	AOI22X1 AOI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5236_), .D(_5255_), .Y(csr_gpr_iu_rs2_9_) );
	NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__10_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5256_) );
	MUX2X1 MUX2X1_97 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__10_), .B(csr_gpr_iu_gpr_29__10_), .S(biu_ins_20_bF_buf0), .Y(_5257_) );
	OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_4911__bF_buf3), .C(_5256_), .Y(_5258_) );
	NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf4), .B(_5258_), .Y(_5259_) );
	NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__10_), .B(_4881__bF_buf11), .Y(_5260_) );
	OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_4899__bF_buf14), .C(_5260_), .Y(_5261_) );
	OAI22X1 OAI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_4896__bF_buf3), .C(_3706_), .D(_4897__bF_buf14), .Y(_5262_) );
	OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_5262_), .B(_5261_), .C(_4903__bF_buf2), .Y(_5263_) );
	NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf3), .B(_5263_), .C(_5259_), .Y(_5264_) );
	OAI22X1 OAI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_4896__bF_buf2), .C(_2817_), .D(_4897__bF_buf13), .Y(_5265_) );
	NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__10_), .B(_4881__bF_buf10), .Y(_5266_) );
	OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_2752_), .B(_4899__bF_buf13), .C(_5266_), .Y(_5267_) );
	OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5267_), .C(_4895__bF_buf3), .Y(_5268_) );
	OAI22X1 OAI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3015_), .B(_4896__bF_buf1), .C(_3715_), .D(_4897__bF_buf12), .Y(_5269_) );
	NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__10_), .B(_4881__bF_buf9), .Y(_5270_) );
	OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_4899__bF_buf12), .C(_5270_), .Y(_5271_) );
	OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(_5271_), .C(_4903__bF_buf1), .Y(_5272_) );
	NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_5268_), .B(_5272_), .C(_4893__bF_buf2), .Y(_5273_) );
	NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5273_), .C(_5264_), .Y(_5274_) );
	OAI22X1 OAI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_4896__bF_buf0), .C(_3683_), .D(_4897__bF_buf11), .Y(_5275_) );
	NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__10_), .B(_4881__bF_buf8), .Y(_5276_) );
	OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_3684_), .B(_4899__bF_buf11), .C(_5276_), .Y(_5277_) );
	OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_5275_), .B(_5277_), .C(_4895__bF_buf2), .Y(_5278_) );
	NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__10_), .B(_4881__bF_buf7), .Y(_5279_) );
	OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .B(_4899__bF_buf10), .C(_5279_), .Y(_5280_) );
	OAI22X1 OAI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_4896__bF_buf13), .C(_3690_), .D(_4897__bF_buf10), .Y(_5281_) );
	OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_5281_), .B(_5280_), .C(_4903__bF_buf0), .Y(_5282_) );
	AOI22X1 AOI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5278_), .D(_5282_), .Y(_5283_) );
	NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__10_), .B(_4881__bF_buf6), .Y(_5284_) );
	OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_4897__bF_buf9), .C(_5284_), .Y(_5285_) );
	OAI22X1 OAI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .B(_4896__bF_buf12), .C(_3672_), .D(_4899__bF_buf9), .Y(_5286_) );
	OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(_5285_), .C(_4895__bF_buf1), .Y(_5287_) );
	NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__10_), .B(_4881__bF_buf5), .Y(_5288_) );
	OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_3678_), .B(_4897__bF_buf8), .C(_5288_), .Y(_5289_) );
	OAI22X1 OAI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(_4896__bF_buf11), .C(_3679_), .D(_4899__bF_buf8), .Y(_5290_) );
	OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5289_), .C(_4903__bF_buf9), .Y(_5291_) );
	AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_5287_), .B(_5291_), .C(_4893__bF_buf1), .Y(_5292_) );
	OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(_5292_), .C(_4931__bF_buf4), .Y(_5293_) );
	AOI22X1 AOI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5274_), .D(_5293_), .Y(csr_gpr_iu_rs2_10_) );
	NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__11_), .B(_4899__bF_buf7), .C(_4897__bF_buf7), .Y(_5294_) );
	MUX2X1 MUX2X1_98 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__11_), .B(csr_gpr_iu_gpr_29__11_), .S(biu_ins_20_bF_buf6), .Y(_5295_) );
	OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_4911__bF_buf2), .C(_5294_), .Y(_5296_) );
	NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf0), .B(_5296_), .Y(_5297_) );
	NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__11_), .B(_4881__bF_buf4), .Y(_5298_) );
	OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_4899__bF_buf6), .C(_5298_), .Y(_5299_) );
	OAI22X1 OAI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_4896__bF_buf10), .C(_3761_), .D(_4897__bF_buf6), .Y(_5300_) );
	OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_5300_), .B(_5299_), .C(_4903__bF_buf8), .Y(_5301_) );
	NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf2), .B(_5301_), .C(_5297_), .Y(_5302_) );
	NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__11_), .B(_4881__bF_buf3), .Y(_5303_) );
	OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .B(_4897__bF_buf5), .C(_5303_), .Y(_5304_) );
	OAI22X1 OAI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_4896__bF_buf9), .C(_2754_), .D(_4899__bF_buf5), .Y(_5305_) );
	OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_5305_), .B(_5304_), .C(_4895__bF_buf10), .Y(_5306_) );
	NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__11_), .B(_4881__bF_buf2), .Y(_5307_) );
	OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_3770_), .B(_4897__bF_buf4), .C(_5307_), .Y(_5308_) );
	OAI22X1 OAI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .B(_4896__bF_buf8), .C(_3771_), .D(_4899__bF_buf4), .Y(_5309_) );
	OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_5309_), .B(_5308_), .C(_4903__bF_buf7), .Y(_5310_) );
	NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_5306_), .B(_5310_), .C(_4893__bF_buf0), .Y(_5311_) );
	NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5311_), .C(_5302_), .Y(_5312_) );
	NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__11_), .B(_4881__bF_buf1), .Y(_5313_) );
	OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .B(_4899__bF_buf3), .C(_5313_), .Y(_5314_) );
	OAI22X1 OAI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_4896__bF_buf7), .C(_3741_), .D(_4897__bF_buf3), .Y(_5315_) );
	OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_5315_), .B(_5314_), .C(_4895__bF_buf9), .Y(_5316_) );
	NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__11_), .B(_4881__bF_buf0), .Y(_5317_) );
	OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_4897__bF_buf2), .C(_5317_), .Y(_5318_) );
	OAI22X1 OAI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .B(_4896__bF_buf6), .C(_3745_), .D(_4899__bF_buf2), .Y(_5319_) );
	OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_5319_), .B(_5318_), .C(_4903__bF_buf6), .Y(_5320_) );
	AOI22X1 AOI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5316_), .D(_5320_), .Y(_5321_) );
	NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__11_), .B(_4881__bF_buf11), .Y(_5322_) );
	OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_4897__bF_buf1), .C(_5322_), .Y(_5323_) );
	OAI22X1 OAI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_4896__bF_buf5), .C(_3727_), .D(_4899__bF_buf1), .Y(_5324_) );
	OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_5324_), .B(_5323_), .C(_4895__bF_buf8), .Y(_5325_) );
	NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__11_), .B(_4881__bF_buf10), .Y(_5326_) );
	OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_3733_), .B(_4897__bF_buf0), .C(_5326_), .Y(_5327_) );
	OAI22X1 OAI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_4896__bF_buf4), .C(_3734_), .D(_4899__bF_buf0), .Y(_5328_) );
	OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_5328_), .B(_5327_), .C(_4903__bF_buf5), .Y(_5329_) );
	AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_5329_), .C(_4893__bF_buf5), .Y(_5330_) );
	OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_5321_), .B(_5330_), .C(_4931__bF_buf3), .Y(_5331_) );
	AOI22X1 AOI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5312_), .D(_5331_), .Y(csr_gpr_iu_rs2_11_) );
	NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__12_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5332_) );
	MUX2X1 MUX2X1_99 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__12_), .B(csr_gpr_iu_gpr_29__12_), .S(biu_ins_20_bF_buf5), .Y(_5333_) );
	OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_5333_), .B(_4911__bF_buf1), .C(_5332_), .Y(_5334_) );
	NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf7), .B(_5334_), .Y(_5335_) );
	NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__12_), .B(_4881__bF_buf9), .Y(_5336_) );
	OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_4899__bF_buf14), .C(_5336_), .Y(_5337_) );
	OAI22X1 OAI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_4896__bF_buf3), .C(_3785_), .D(_4897__bF_buf14), .Y(_5338_) );
	OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_5338_), .B(_5337_), .C(_4903__bF_buf4), .Y(_5339_) );
	NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf1), .B(_5339_), .C(_5335_), .Y(_5340_) );
	OAI22X1 OAI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .B(_4896__bF_buf2), .C(_2821_), .D(_4897__bF_buf13), .Y(_5341_) );
	NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__12_), .B(_4881__bF_buf8), .Y(_5342_) );
	OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_4899__bF_buf13), .C(_5342_), .Y(_5343_) );
	OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_5341_), .B(_5343_), .C(_4895__bF_buf6), .Y(_5344_) );
	OAI22X1 OAI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_4896__bF_buf1), .C(_3794_), .D(_4897__bF_buf12), .Y(_5345_) );
	NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__12_), .B(_4881__bF_buf7), .Y(_5346_) );
	OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_4899__bF_buf12), .C(_5346_), .Y(_5347_) );
	OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_5345_), .B(_5347_), .C(_4903__bF_buf3), .Y(_5348_) );
	NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_5344_), .B(_5348_), .C(_4893__bF_buf4), .Y(_5349_) );
	NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5349_), .C(_5340_), .Y(_5350_) );
	NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__12_), .B(_4881__bF_buf6), .Y(_5351_) );
	OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_3802_), .B(_4897__bF_buf11), .C(_5351_), .Y(_5352_) );
	OAI22X1 OAI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(_4896__bF_buf0), .C(_3805_), .D(_4899__bF_buf11), .Y(_5353_) );
	OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_5352_), .C(_4895__bF_buf5), .Y(_5354_) );
	NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__12_), .B(_4881__bF_buf5), .Y(_5355_) );
	OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_3809_), .B(_4899__bF_buf10), .C(_5355_), .Y(_5356_) );
	OAI22X1 OAI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_4896__bF_buf13), .C(_3812_), .D(_4897__bF_buf10), .Y(_5357_) );
	OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_5357_), .B(_5356_), .C(_4903__bF_buf2), .Y(_5358_) );
	AOI22X1 AOI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5354_), .D(_5358_), .Y(_5359_) );
	NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__12_), .B(_4881__bF_buf4), .Y(_5360_) );
	OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(_4897__bF_buf9), .C(_5360_), .Y(_5361_) );
	OAI22X1 OAI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_4896__bF_buf12), .C(_3820_), .D(_4899__bF_buf9), .Y(_5362_) );
	OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_5362_), .B(_5361_), .C(_4895__bF_buf4), .Y(_5363_) );
	NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__12_), .B(_4881__bF_buf3), .Y(_5364_) );
	OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_4897__bF_buf8), .C(_5364_), .Y(_5365_) );
	OAI22X1 OAI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_4896__bF_buf11), .C(_3827_), .D(_4899__bF_buf8), .Y(_5366_) );
	OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_5366_), .B(_5365_), .C(_4903__bF_buf1), .Y(_5367_) );
	AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_5367_), .C(_4893__bF_buf3), .Y(_5368_) );
	OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_5359_), .B(_5368_), .C(_4931__bF_buf2), .Y(_5369_) );
	AOI22X1 AOI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5350_), .D(_5369_), .Y(csr_gpr_iu_rs2_12_) );
	OAI22X1 OAI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(_4896__bF_buf10), .C(_3833_), .D(_4891__bF_buf1), .Y(_5370_) );
	OAI22X1 OAI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_4897__bF_buf7), .C(_3837_), .D(_4899__bF_buf7), .Y(_5371_) );
	OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_5370_), .B(_5371_), .C(_4895__bF_buf3), .Y(_5372_) );
	OAI22X1 OAI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_4896__bF_buf9), .C(_3840_), .D(_4891__bF_buf0), .Y(_5373_) );
	OAI22X1 OAI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_4897__bF_buf6), .C(_3844_), .D(_4899__bF_buf6), .Y(_5374_) );
	OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_5373_), .B(_5374_), .C(_4903__bF_buf0), .Y(_5375_) );
	AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5372_), .C(_4893__bF_buf2), .Y(_5376_) );
	NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__13_), .B(_4881__bF_buf2), .Y(_5377_) );
	OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .B(_4899__bF_buf5), .C(_5377_), .Y(_5378_) );
	OAI22X1 OAI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_4896__bF_buf8), .C(_3851_), .D(_4897__bF_buf5), .Y(_5379_) );
	OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_5379_), .B(_5378_), .C(_4895__bF_buf2), .Y(_5380_) );
	NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__13_), .B(_4881__bF_buf1), .Y(_5381_) );
	OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .B(_4899__bF_buf4), .C(_5381_), .Y(_5382_) );
	OAI22X1 OAI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(_4896__bF_buf7), .C(_3858_), .D(_4897__bF_buf4), .Y(_5383_) );
	OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_5382_), .C(_4903__bF_buf9), .Y(_5384_) );
	AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .B(_5384_), .C(_4910__bF_buf0), .Y(_5385_) );
	OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_5376_), .B(_5385_), .C(_4931__bF_buf1), .Y(_5386_) );
	OAI22X1 OAI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .B(_4897__bF_buf3), .C(_3865_), .D(_4899__bF_buf3), .Y(_5387_) );
	NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__13_), .B(biu_ins_20_bF_buf4), .Y(_5388_) );
	OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(_3867_), .C(_5388_), .Y(_5389_) );
	AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf0), .B(_5389_), .C(_5387_), .Y(_5390_) );
	OAI22X1 OAI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_4897__bF_buf2), .C(_3872_), .D(_4899__bF_buf2), .Y(_5391_) );
	AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__13_), .B(_4911__bF_buf5), .C(_5391_), .Y(_5392_) );
	MUX2X1 MUX2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_5392_), .B(_5390_), .S(_4895__bF_buf1), .Y(_5393_) );
	NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__13_), .B(_4881__bF_buf0), .Y(_5394_) );
	OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_4897__bF_buf1), .C(_5394_), .Y(_5395_) );
	OAI22X1 OAI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_4896__bF_buf6), .C(_2758_), .D(_4899__bF_buf1), .Y(_5396_) );
	OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_5396_), .B(_5395_), .C(_4895__bF_buf0), .Y(_5397_) );
	OAI22X1 OAI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3880_), .B(_4897__bF_buf0), .C(_3881_), .D(_4899__bF_buf0), .Y(_5398_) );
	OAI22X1 OAI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_4896__bF_buf5), .C(_3883_), .D(_4891__bF_buf7), .Y(_5399_) );
	OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_5399_), .B(_5398_), .C(_4903__bF_buf8), .Y(_5400_) );
	AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_5397_), .B(_5400_), .C(_4910__bF_buf7), .Y(_5401_) );
	AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .B(_4910__bF_buf6), .C(_5401_), .Y(_5402_) );
	OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf1), .B(_5402_), .C(_5386_), .Y(csr_gpr_iu_rs2_13_) );
	OAI22X1 OAI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_4896__bF_buf4), .C(_3888_), .D(_4891__bF_buf6), .Y(_5403_) );
	OAI22X1 OAI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_4897__bF_buf15), .C(_3892_), .D(_4899__bF_buf15), .Y(_5404_) );
	OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .B(_5404_), .C(_4895__bF_buf10), .Y(_5405_) );
	OAI22X1 OAI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3896_), .B(_4896__bF_buf3), .C(_3895_), .D(_4891__bF_buf5), .Y(_5406_) );
	OAI22X1 OAI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(_4897__bF_buf14), .C(_3899_), .D(_4899__bF_buf14), .Y(_5407_) );
	OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .B(_5407_), .C(_4903__bF_buf7), .Y(_5408_) );
	AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .B(_5405_), .C(_4893__bF_buf1), .Y(_5409_) );
	NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__14_), .B(_4881__bF_buf11), .Y(_5410_) );
	OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(_4899__bF_buf13), .C(_5410_), .Y(_5411_) );
	OAI22X1 OAI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3904_), .B(_4896__bF_buf2), .C(_3906_), .D(_4897__bF_buf13), .Y(_5412_) );
	OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_5412_), .B(_5411_), .C(_4895__bF_buf9), .Y(_5413_) );
	NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__14_), .B(_4881__bF_buf10), .Y(_5414_) );
	OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_3910_), .B(_4899__bF_buf12), .C(_5414_), .Y(_5415_) );
	OAI22X1 OAI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_4896__bF_buf1), .C(_3913_), .D(_4897__bF_buf12), .Y(_5416_) );
	OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_5416_), .B(_5415_), .C(_4903__bF_buf6), .Y(_5417_) );
	AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_5413_), .B(_5417_), .C(_4910__bF_buf5), .Y(_5418_) );
	OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_5409_), .B(_5418_), .C(_4931__bF_buf0), .Y(_5419_) );
	OAI22X1 OAI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_4897__bF_buf11), .C(_3920_), .D(_4899__bF_buf11), .Y(_5420_) );
	NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__14_), .B(biu_ins_20_bF_buf2), .Y(_5421_) );
	OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf1), .B(_3922_), .C(_5421_), .Y(_5422_) );
	AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf4), .B(_5422_), .C(_5420_), .Y(_5423_) );
	OAI22X1 OAI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_4897__bF_buf10), .C(_3927_), .D(_4899__bF_buf10), .Y(_5424_) );
	AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__14_), .B(_4911__bF_buf3), .C(_5424_), .Y(_5425_) );
	MUX2X1 MUX2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .B(_5423_), .S(_4895__bF_buf8), .Y(_5426_) );
	OAI22X1 OAI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_4896__bF_buf0), .C(_2825_), .D(_4897__bF_buf9), .Y(_5427_) );
	NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__14_), .B(_4881__bF_buf9), .Y(_5428_) );
	OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_4899__bF_buf9), .C(_5428_), .Y(_5429_) );
	OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_5429_), .C(_4895__bF_buf7), .Y(_5430_) );
	OAI22X1 OAI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_4897__bF_buf8), .C(_3936_), .D(_4899__bF_buf8), .Y(_5431_) );
	OAI22X1 OAI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_4896__bF_buf13), .C(_3938_), .D(_4891__bF_buf4), .Y(_5432_) );
	OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_5432_), .B(_5431_), .C(_4903__bF_buf5), .Y(_5433_) );
	AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_5430_), .B(_5433_), .C(_4910__bF_buf4), .Y(_5434_) );
	AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_5426_), .B(_4910__bF_buf3), .C(_5434_), .Y(_5435_) );
	OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf0), .B(_5435_), .C(_5419_), .Y(csr_gpr_iu_rs2_14_) );
	OAI22X1 OAI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3944_), .B(_4896__bF_buf12), .C(_3943_), .D(_4891__bF_buf3), .Y(_5436_) );
	OAI22X1 OAI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_4897__bF_buf7), .C(_3947_), .D(_4899__bF_buf7), .Y(_5437_) );
	OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_5436_), .B(_5437_), .C(_4895__bF_buf6), .Y(_5438_) );
	OAI22X1 OAI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_4896__bF_buf11), .C(_3950_), .D(_4891__bF_buf2), .Y(_5439_) );
	OAI22X1 OAI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_4897__bF_buf6), .C(_3954_), .D(_4899__bF_buf6), .Y(_5440_) );
	OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_5439_), .B(_5440_), .C(_4903__bF_buf4), .Y(_5441_) );
	AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_5441_), .B(_5438_), .C(_4893__bF_buf0), .Y(_5442_) );
	OAI22X1 OAI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_4896__bF_buf10), .C(_3958_), .D(_4899__bF_buf5), .Y(_5443_) );
	NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__15_), .B(_4881__bF_buf8), .Y(_5444_) );
	OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_4897__bF_buf5), .C(_5444_), .Y(_5445_) );
	OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_5445_), .C(_4895__bF_buf5), .Y(_5446_) );
	OAI22X1 OAI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3966_), .B(_4896__bF_buf9), .C(_3965_), .D(_4899__bF_buf4), .Y(_5447_) );
	NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__15_), .B(_4881__bF_buf7), .Y(_5448_) );
	OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_4897__bF_buf4), .C(_5448_), .Y(_5449_) );
	OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_5447_), .B(_5449_), .C(_4903__bF_buf3), .Y(_5450_) );
	AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_5446_), .B(_5450_), .C(_4910__bF_buf2), .Y(_5451_) );
	OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_5442_), .B(_5451_), .C(_4931__bF_buf4), .Y(_5452_) );
	OAI22X1 OAI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3974_), .B(_4897__bF_buf3), .C(_3975_), .D(_4899__bF_buf3), .Y(_5453_) );
	NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__15_), .B(biu_ins_20_bF_buf0), .Y(_5454_) );
	OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf6), .B(_3977_), .C(_5454_), .Y(_5455_) );
	AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf2), .B(_5455_), .C(_5453_), .Y(_5456_) );
	OAI22X1 OAI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3981_), .B(_4897__bF_buf2), .C(_3982_), .D(_4899__bF_buf2), .Y(_5457_) );
	AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__15_), .B(_4911__bF_buf1), .C(_5457_), .Y(_5458_) );
	MUX2X1 MUX2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_5458_), .B(_5456_), .S(_4895__bF_buf4), .Y(_5459_) );
	OAI22X1 OAI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2892_), .B(_4896__bF_buf8), .C(_2827_), .D(_4897__bF_buf1), .Y(_5460_) );
	NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__15_), .B(_4881__bF_buf6), .Y(_5461_) );
	OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_4899__bF_buf1), .C(_5461_), .Y(_5462_) );
	OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_5460_), .B(_5462_), .C(_4895__bF_buf3), .Y(_5463_) );
	OAI22X1 OAI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_4897__bF_buf0), .C(_3991_), .D(_4899__bF_buf0), .Y(_5464_) );
	OAI22X1 OAI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_4896__bF_buf7), .C(_3993_), .D(_4891__bF_buf1), .Y(_5465_) );
	OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_5465_), .B(_5464_), .C(_4903__bF_buf2), .Y(_5466_) );
	AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_5463_), .B(_5466_), .C(_4910__bF_buf1), .Y(_5467_) );
	AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_5459_), .B(_4910__bF_buf0), .C(_5467_), .Y(_5468_) );
	OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf3), .B(_5468_), .C(_5452_), .Y(csr_gpr_iu_rs2_15_) );
	NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__16_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5469_) );
	MUX2X1 MUX2X1_103 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__16_), .B(csr_gpr_iu_gpr_29__16_), .S(biu_ins_20_bF_buf5), .Y(_5470_) );
	OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_5470_), .B(_4911__bF_buf0), .C(_5469_), .Y(_5471_) );
	NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf2), .B(_5471_), .Y(_5472_) );
	NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__16_), .B(_4881__bF_buf5), .Y(_5473_) );
	OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_4002_), .B(_4899__bF_buf14), .C(_5473_), .Y(_5474_) );
	OAI22X1 OAI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_4896__bF_buf6), .C(_4005_), .D(_4897__bF_buf14), .Y(_5475_) );
	OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_5475_), .B(_5474_), .C(_4903__bF_buf1), .Y(_5476_) );
	NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_5476_), .C(_5472_), .Y(_5477_) );
	NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__16_), .B(_4881__bF_buf4), .Y(_5478_) );
	OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_2829_), .B(_4897__bF_buf13), .C(_5478_), .Y(_5479_) );
	OAI22X1 OAI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_4896__bF_buf5), .C(_2764_), .D(_4899__bF_buf13), .Y(_5480_) );
	OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_5480_), .B(_5479_), .C(_4895__bF_buf1), .Y(_5481_) );
	NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__16_), .B(_4881__bF_buf3), .Y(_5482_) );
	OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_4897__bF_buf12), .C(_5482_), .Y(_5483_) );
	OAI22X1 OAI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_4896__bF_buf4), .C(_4016_), .D(_4899__bF_buf12), .Y(_5484_) );
	OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_5484_), .B(_5483_), .C(_4903__bF_buf0), .Y(_5485_) );
	NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_5481_), .B(_5485_), .C(_4893__bF_buf5), .Y(_5486_) );
	NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5486_), .C(_5477_), .Y(_5487_) );
	NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__16_), .B(_4881__bF_buf2), .Y(_5488_) );
	OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_4897__bF_buf11), .C(_5488_), .Y(_5489_) );
	OAI22X1 OAI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .B(_4896__bF_buf3), .C(_4025_), .D(_4899__bF_buf11), .Y(_5490_) );
	OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_5490_), .B(_5489_), .C(_4895__bF_buf0), .Y(_5491_) );
	NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__16_), .B(_4881__bF_buf1), .Y(_5492_) );
	OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_4029_), .B(_4899__bF_buf10), .C(_5492_), .Y(_5493_) );
	OAI22X1 OAI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .B(_4896__bF_buf2), .C(_4032_), .D(_4897__bF_buf10), .Y(_5494_) );
	OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_5494_), .B(_5493_), .C(_4903__bF_buf9), .Y(_5495_) );
	AOI22X1 AOI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5491_), .D(_5495_), .Y(_5496_) );
	NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__16_), .B(_4881__bF_buf0), .Y(_5497_) );
	OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(_4897__bF_buf9), .C(_5497_), .Y(_5498_) );
	OAI22X1 OAI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(_4041_), .B(_4896__bF_buf1), .C(_4040_), .D(_4899__bF_buf9), .Y(_5499_) );
	OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .B(_5498_), .C(_4895__bF_buf10), .Y(_5500_) );
	NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__16_), .B(_4881__bF_buf11), .Y(_5501_) );
	OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_4044_), .B(_4897__bF_buf8), .C(_5501_), .Y(_5502_) );
	OAI22X1 OAI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_4896__bF_buf0), .C(_4047_), .D(_4899__bF_buf8), .Y(_5503_) );
	OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5502_), .C(_4903__bF_buf8), .Y(_5504_) );
	AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_5500_), .B(_5504_), .C(_4893__bF_buf4), .Y(_5505_) );
	OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_5496_), .B(_5505_), .C(_4931__bF_buf3), .Y(_5506_) );
	AOI22X1 AOI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5487_), .D(_5506_), .Y(csr_gpr_iu_rs2_16_) );
	NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__17_), .B(_4899__bF_buf7), .C(_4897__bF_buf7), .Y(_5507_) );
	MUX2X1 MUX2X1_104 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__17_), .B(csr_gpr_iu_gpr_29__17_), .S(biu_ins_20_bF_buf4), .Y(_5508_) );
	OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_4911__bF_buf5), .C(_5507_), .Y(_5509_) );
	NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf9), .B(_5509_), .Y(_5510_) );
	NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__17_), .B(_4881__bF_buf10), .Y(_5511_) );
	OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .B(_4899__bF_buf6), .C(_5511_), .Y(_5512_) );
	OAI22X1 OAI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(_4061_), .B(_4896__bF_buf13), .C(_4060_), .D(_4897__bF_buf6), .Y(_5513_) );
	OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_5513_), .B(_5512_), .C(_4903__bF_buf7), .Y(_5514_) );
	NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf6), .B(_5514_), .C(_5510_), .Y(_5515_) );
	NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__17_), .B(_4881__bF_buf9), .Y(_5516_) );
	OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_4897__bF_buf5), .C(_5516_), .Y(_5517_) );
	OAI22X1 OAI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_4896__bF_buf12), .C(_2766_), .D(_4899__bF_buf5), .Y(_5518_) );
	OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_5518_), .B(_5517_), .C(_4895__bF_buf8), .Y(_5519_) );
	NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__17_), .B(_4881__bF_buf8), .Y(_5520_) );
	OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_4897__bF_buf4), .C(_5520_), .Y(_5521_) );
	OAI22X1 OAI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .B(_4896__bF_buf11), .C(_4072_), .D(_4899__bF_buf4), .Y(_5522_) );
	OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_5522_), .B(_5521_), .C(_4903__bF_buf6), .Y(_5523_) );
	NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_5519_), .B(_5523_), .C(_4893__bF_buf3), .Y(_5524_) );
	NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5524_), .C(_5515_), .Y(_5525_) );
	NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__17_), .B(_4881__bF_buf7), .Y(_5526_) );
	OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_4077_), .B(_4897__bF_buf3), .C(_5526_), .Y(_5527_) );
	OAI22X1 OAI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(_4896__bF_buf10), .C(_4080_), .D(_4899__bF_buf3), .Y(_5528_) );
	OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_5528_), .B(_5527_), .C(_4895__bF_buf7), .Y(_5529_) );
	NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__17_), .B(_4881__bF_buf6), .Y(_5530_) );
	OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .B(_4899__bF_buf2), .C(_5530_), .Y(_5531_) );
	OAI22X1 OAI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .B(_4896__bF_buf9), .C(_4087_), .D(_4897__bF_buf2), .Y(_5532_) );
	OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_5532_), .B(_5531_), .C(_4903__bF_buf5), .Y(_5533_) );
	AOI22X1 AOI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5529_), .D(_5533_), .Y(_5534_) );
	NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__17_), .B(_4881__bF_buf5), .Y(_5535_) );
	OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_4092_), .B(_4897__bF_buf1), .C(_5535_), .Y(_5536_) );
	OAI22X1 OAI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_4896__bF_buf8), .C(_4095_), .D(_4899__bF_buf1), .Y(_5537_) );
	OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_5537_), .B(_5536_), .C(_4895__bF_buf6), .Y(_5538_) );
	NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__17_), .B(_4881__bF_buf4), .Y(_5539_) );
	OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_4897__bF_buf0), .C(_5539_), .Y(_5540_) );
	OAI22X1 OAI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .B(_4896__bF_buf7), .C(_4102_), .D(_4899__bF_buf0), .Y(_5541_) );
	OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_5541_), .B(_5540_), .C(_4903__bF_buf4), .Y(_5542_) );
	AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_5538_), .B(_5542_), .C(_4893__bF_buf2), .Y(_5543_) );
	OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_5534_), .B(_5543_), .C(_4931__bF_buf2), .Y(_5544_) );
	AOI22X1 AOI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5525_), .D(_5544_), .Y(csr_gpr_iu_rs2_17_) );
	OAI22X1 OAI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_4896__bF_buf6), .C(_4151_), .D(_4891__bF_buf0), .Y(_5545_) );
	OAI22X1 OAI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(_4147_), .B(_4897__bF_buf15), .C(_4150_), .D(_4899__bF_buf15), .Y(_5546_) );
	OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_5545_), .B(_5546_), .C(_4895__bF_buf5), .Y(_5547_) );
	OAI22X1 OAI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4896__bF_buf5), .C(_4158_), .D(_4891__bF_buf7), .Y(_5548_) );
	OAI22X1 OAI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(_4154_), .B(_4897__bF_buf14), .C(_4157_), .D(_4899__bF_buf14), .Y(_5549_) );
	OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_5548_), .B(_5549_), .C(_4903__bF_buf3), .Y(_5550_) );
	AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_5550_), .B(_5547_), .C(_4893__bF_buf1), .Y(_5551_) );
	NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__18_), .B(_4881__bF_buf3), .Y(_5552_) );
	OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .B(_4899__bF_buf13), .C(_5552_), .Y(_5553_) );
	OAI22X1 OAI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_4896__bF_buf4), .C(_4132_), .D(_4897__bF_buf13), .Y(_5554_) );
	OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_5554_), .B(_5553_), .C(_4895__bF_buf4), .Y(_5555_) );
	NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__18_), .B(_4881__bF_buf2), .Y(_5556_) );
	OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_4899__bF_buf12), .C(_5556_), .Y(_5557_) );
	OAI22X1 OAI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(_4143_), .B(_4896__bF_buf3), .C(_4142_), .D(_4897__bF_buf12), .Y(_5558_) );
	OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_5558_), .B(_5557_), .C(_4903__bF_buf2), .Y(_5559_) );
	AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_5555_), .B(_5559_), .C(_4910__bF_buf5), .Y(_5560_) );
	OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_5560_), .C(_4931__bF_buf1), .Y(_5561_) );
	INVX1 INVX1_1109 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__18_), .Y(_5562_) );
	INVX1 INVX1_1110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__18_), .Y(_5563_) );
	OAI22X1 OAI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(_5562_), .B(_4897__bF_buf11), .C(_5563_), .D(_4899__bF_buf11), .Y(_5564_) );
	AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__18_), .B(_4911__bF_buf4), .C(_5564_), .Y(_5565_) );
	OAI22X1 OAI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .B(_4899__bF_buf10), .C(_4112_), .D(_4891__bF_buf6), .Y(_5566_) );
	OAI22X1 OAI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .B(_4896__bF_buf2), .C(_4115_), .D(_4897__bF_buf10), .Y(_5567_) );
	OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_5566_), .B(_5567_), .C(_4903__bF_buf1), .Y(_5568_) );
	OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_4903__bF_buf0), .B(_5565_), .C(_5568_), .Y(_5569_) );
	OAI22X1 OAI22X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_4896__bF_buf1), .C(_2833_), .D(_4897__bF_buf9), .Y(_5570_) );
	NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__18_), .B(_4881__bF_buf1), .Y(_5571_) );
	OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_4899__bF_buf9), .C(_5571_), .Y(_5572_) );
	OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_5570_), .B(_5572_), .C(_4895__bF_buf3), .Y(_5573_) );
	OAI22X1 OAI22X1_507 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(_4897__bF_buf8), .C(_4127_), .D(_4899__bF_buf8), .Y(_5574_) );
	OAI22X1 OAI22X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_4896__bF_buf0), .C(_4126_), .D(_4891__bF_buf5), .Y(_5575_) );
	OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_5575_), .B(_5574_), .C(_4903__bF_buf9), .Y(_5576_) );
	AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_5576_), .C(_4910__bF_buf4), .Y(_5577_) );
	AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_5569_), .B(_4910__bF_buf3), .C(_5577_), .Y(_5578_) );
	OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf2), .B(_5578_), .C(_5561_), .Y(csr_gpr_iu_rs2_18_) );
	OAI22X1 OAI22X1_509 ( .gnd(gnd), .vdd(vdd), .A(_4164_), .B(_4896__bF_buf13), .C(_4163_), .D(_4891__bF_buf4), .Y(_5579_) );
	OAI22X1 OAI22X1_510 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_4897__bF_buf7), .C(_4167_), .D(_4899__bF_buf7), .Y(_5580_) );
	OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_5579_), .B(_5580_), .C(_4895__bF_buf2), .Y(_5581_) );
	OAI22X1 OAI22X1_511 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .B(_4896__bF_buf12), .C(_4170_), .D(_4891__bF_buf3), .Y(_5582_) );
	OAI22X1 OAI22X1_512 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_4897__bF_buf6), .C(_4174_), .D(_4899__bF_buf6), .Y(_5583_) );
	OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_5582_), .B(_5583_), .C(_4903__bF_buf8), .Y(_5584_) );
	AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_5584_), .B(_5581_), .C(_4893__bF_buf0), .Y(_5585_) );
	OAI22X1 OAI22X1_513 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .B(_4896__bF_buf11), .C(_4178_), .D(_4899__bF_buf5), .Y(_5586_) );
	NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__19_), .B(_4881__bF_buf0), .Y(_5587_) );
	OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_4181_), .B(_4897__bF_buf5), .C(_5587_), .Y(_5588_) );
	OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_5586_), .B(_5588_), .C(_4895__bF_buf1), .Y(_5589_) );
	OAI22X1 OAI22X1_514 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .B(_4896__bF_buf10), .C(_4185_), .D(_4899__bF_buf4), .Y(_5590_) );
	NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__19_), .B(_4881__bF_buf11), .Y(_5591_) );
	OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_4188_), .B(_4897__bF_buf4), .C(_5591_), .Y(_5592_) );
	OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_5590_), .B(_5592_), .C(_4903__bF_buf7), .Y(_5593_) );
	AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_5589_), .B(_5593_), .C(_4910__bF_buf2), .Y(_5594_) );
	OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_5585_), .B(_5594_), .C(_4931__bF_buf0), .Y(_5595_) );
	OAI22X1 OAI22X1_515 ( .gnd(gnd), .vdd(vdd), .A(_4194_), .B(_4897__bF_buf3), .C(_4195_), .D(_4899__bF_buf3), .Y(_5596_) );
	NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__19_), .B(biu_ins_20_bF_buf3), .Y(_5597_) );
	OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf2), .B(_4197_), .C(_5597_), .Y(_5598_) );
	AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf3), .B(_5598_), .C(_5596_), .Y(_5599_) );
	OAI22X1 OAI22X1_516 ( .gnd(gnd), .vdd(vdd), .A(_4201_), .B(_4897__bF_buf2), .C(_4202_), .D(_4899__bF_buf2), .Y(_5600_) );
	AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__19_), .B(_4911__bF_buf2), .C(_5600_), .Y(_5601_) );
	MUX2X1 MUX2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_5601_), .B(_5599_), .S(_4895__bF_buf0), .Y(_5602_) );
	OAI22X1 OAI22X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_4896__bF_buf9), .C(_2835_), .D(_4897__bF_buf1), .Y(_5603_) );
	NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__19_), .B(_4881__bF_buf10), .Y(_5604_) );
	OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_2770_), .B(_4899__bF_buf1), .C(_5604_), .Y(_5605_) );
	OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_5603_), .B(_5605_), .C(_4895__bF_buf10), .Y(_5606_) );
	OAI22X1 OAI22X1_518 ( .gnd(gnd), .vdd(vdd), .A(_4210_), .B(_4897__bF_buf0), .C(_4211_), .D(_4899__bF_buf0), .Y(_5607_) );
	OAI22X1 OAI22X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .B(_4896__bF_buf8), .C(_4213_), .D(_4891__bF_buf2), .Y(_5608_) );
	OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_5608_), .B(_5607_), .C(_4903__bF_buf6), .Y(_5609_) );
	AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_5606_), .B(_5609_), .C(_4910__bF_buf1), .Y(_5610_) );
	AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_5602_), .B(_4910__bF_buf0), .C(_5610_), .Y(_5611_) );
	OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf1), .B(_5611_), .C(_5595_), .Y(csr_gpr_iu_rs2_19_) );
	NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__20_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5612_) );
	MUX2X1 MUX2X1_106 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__20_), .B(csr_gpr_iu_gpr_29__20_), .S(biu_ins_20_bF_buf1), .Y(_5613_) );
	OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .B(_4911__bF_buf1), .C(_5612_), .Y(_5614_) );
	NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf9), .B(_5614_), .Y(_5615_) );
	NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__20_), .B(_4881__bF_buf9), .Y(_5616_) );
	OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_4222_), .B(_4899__bF_buf14), .C(_5616_), .Y(_5617_) );
	OAI22X1 OAI22X1_520 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4896__bF_buf7), .C(_4225_), .D(_4897__bF_buf14), .Y(_5618_) );
	OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_5618_), .B(_5617_), .C(_4903__bF_buf5), .Y(_5619_) );
	NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_5619_), .C(_5615_), .Y(_5620_) );
	OAI22X1 OAI22X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_4896__bF_buf6), .C(_2837_), .D(_4897__bF_buf13), .Y(_5621_) );
	NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__20_), .B(_4881__bF_buf8), .Y(_5622_) );
	OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_4899__bF_buf13), .C(_5622_), .Y(_5623_) );
	OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_5621_), .B(_5623_), .C(_4895__bF_buf8), .Y(_5624_) );
	OAI22X1 OAI22X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_4896__bF_buf5), .C(_4234_), .D(_4897__bF_buf12), .Y(_5625_) );
	NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__20_), .B(_4881__bF_buf7), .Y(_5626_) );
	OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_4899__bF_buf12), .C(_5626_), .Y(_5627_) );
	OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_5625_), .B(_5627_), .C(_4903__bF_buf4), .Y(_5628_) );
	NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_5624_), .B(_5628_), .C(_4893__bF_buf5), .Y(_5629_) );
	NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5629_), .C(_5620_), .Y(_5630_) );
	OAI22X1 OAI22X1_523 ( .gnd(gnd), .vdd(vdd), .A(_4246_), .B(_4896__bF_buf4), .C(_4242_), .D(_4897__bF_buf11), .Y(_5631_) );
	NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__20_), .B(_4881__bF_buf6), .Y(_5632_) );
	OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_4245_), .B(_4899__bF_buf11), .C(_5632_), .Y(_5633_) );
	OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_5631_), .B(_5633_), .C(_4895__bF_buf7), .Y(_5634_) );
	OAI22X1 OAI22X1_524 ( .gnd(gnd), .vdd(vdd), .A(_4250_), .B(_4896__bF_buf3), .C(_4249_), .D(_4899__bF_buf10), .Y(_5635_) );
	NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__20_), .B(_4881__bF_buf5), .Y(_5636_) );
	OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_4252_), .B(_4897__bF_buf10), .C(_5636_), .Y(_5637_) );
	OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_5637_), .C(_4903__bF_buf3), .Y(_5638_) );
	AOI22X1 AOI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5634_), .D(_5638_), .Y(_5639_) );
	OAI22X1 OAI22X1_525 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(_4896__bF_buf2), .C(_4257_), .D(_4897__bF_buf9), .Y(_5640_) );
	NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__20_), .B(_4881__bF_buf4), .Y(_5641_) );
	OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_4260_), .B(_4899__bF_buf9), .C(_5641_), .Y(_5642_) );
	OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_5640_), .B(_5642_), .C(_4895__bF_buf6), .Y(_5643_) );
	OAI22X1 OAI22X1_526 ( .gnd(gnd), .vdd(vdd), .A(_4268_), .B(_4896__bF_buf1), .C(_4264_), .D(_4897__bF_buf8), .Y(_5644_) );
	NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__20_), .B(_4881__bF_buf3), .Y(_5645_) );
	OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_4267_), .B(_4899__bF_buf8), .C(_5645_), .Y(_5646_) );
	OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_5644_), .B(_5646_), .C(_4903__bF_buf2), .Y(_5647_) );
	AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_5643_), .B(_5647_), .C(_4893__bF_buf4), .Y(_5648_) );
	OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_5639_), .B(_5648_), .C(_4931__bF_buf4), .Y(_5649_) );
	AOI22X1 AOI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5630_), .D(_5649_), .Y(csr_gpr_iu_rs2_20_) );
	OAI22X1 OAI22X1_527 ( .gnd(gnd), .vdd(vdd), .A(_4274_), .B(_4896__bF_buf0), .C(_4273_), .D(_4891__bF_buf1), .Y(_5650_) );
	OAI22X1 OAI22X1_528 ( .gnd(gnd), .vdd(vdd), .A(_4276_), .B(_4897__bF_buf7), .C(_4277_), .D(_4899__bF_buf7), .Y(_5651_) );
	OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_5650_), .B(_5651_), .C(_4895__bF_buf5), .Y(_5652_) );
	OAI22X1 OAI22X1_529 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_4896__bF_buf13), .C(_4280_), .D(_4891__bF_buf0), .Y(_5653_) );
	OAI22X1 OAI22X1_530 ( .gnd(gnd), .vdd(vdd), .A(_4283_), .B(_4897__bF_buf6), .C(_4284_), .D(_4899__bF_buf6), .Y(_5654_) );
	OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_5654_), .C(_4903__bF_buf1), .Y(_5655_) );
	AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_5655_), .B(_5652_), .C(_4893__bF_buf3), .Y(_5656_) );
	OAI22X1 OAI22X1_531 ( .gnd(gnd), .vdd(vdd), .A(_4288_), .B(_4897__bF_buf5), .C(_4289_), .D(_4899__bF_buf5), .Y(_5657_) );
	OAI22X1 OAI22X1_532 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .B(_4896__bF_buf12), .C(_4291_), .D(_4891__bF_buf7), .Y(_5658_) );
	OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_5658_), .B(_5657_), .C(_4895__bF_buf4), .Y(_5659_) );
	OAI22X1 OAI22X1_533 ( .gnd(gnd), .vdd(vdd), .A(_4295_), .B(_4897__bF_buf4), .C(_4296_), .D(_4899__bF_buf4), .Y(_5660_) );
	OAI22X1 OAI22X1_534 ( .gnd(gnd), .vdd(vdd), .A(_4299_), .B(_4896__bF_buf11), .C(_4298_), .D(_4891__bF_buf6), .Y(_5661_) );
	OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_5661_), .B(_5660_), .C(_4903__bF_buf0), .Y(_5662_) );
	AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_5662_), .B(_5659_), .C(_4910__bF_buf6), .Y(_5663_) );
	OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_5656_), .B(_5663_), .C(_4931__bF_buf3), .Y(_5664_) );
	OAI22X1 OAI22X1_535 ( .gnd(gnd), .vdd(vdd), .A(_4304_), .B(_4897__bF_buf3), .C(_4305_), .D(_4899__bF_buf3), .Y(_5665_) );
	NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__21_), .B(biu_ins_20_bF_buf0), .Y(_5666_) );
	OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf6), .B(_4307_), .C(_5666_), .Y(_5667_) );
	AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf0), .B(_5667_), .C(_5665_), .Y(_5668_) );
	OAI22X1 OAI22X1_536 ( .gnd(gnd), .vdd(vdd), .A(_4311_), .B(_4897__bF_buf2), .C(_4312_), .D(_4899__bF_buf2), .Y(_5669_) );
	AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__21_), .B(_4911__bF_buf5), .C(_5669_), .Y(_5670_) );
	MUX2X1 MUX2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_5670_), .B(_5668_), .S(_4895__bF_buf3), .Y(_5671_) );
	NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__21_), .B(_4881__bF_buf2), .Y(_5672_) );
	OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_4897__bF_buf1), .C(_5672_), .Y(_5673_) );
	OAI22X1 OAI22X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(_4896__bF_buf10), .C(_2774_), .D(_4899__bF_buf1), .Y(_5674_) );
	OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_5674_), .B(_5673_), .C(_4895__bF_buf2), .Y(_5675_) );
	OAI22X1 OAI22X1_538 ( .gnd(gnd), .vdd(vdd), .A(_4320_), .B(_4897__bF_buf0), .C(_4321_), .D(_4899__bF_buf0), .Y(_5676_) );
	OAI22X1 OAI22X1_539 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_4896__bF_buf9), .C(_4323_), .D(_4891__bF_buf5), .Y(_5677_) );
	OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_5677_), .B(_5676_), .C(_4903__bF_buf9), .Y(_5678_) );
	AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_5675_), .B(_5678_), .C(_4910__bF_buf5), .Y(_5679_) );
	AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_5671_), .B(_4910__bF_buf4), .C(_5679_), .Y(_5680_) );
	OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf0), .B(_5680_), .C(_5664_), .Y(csr_gpr_iu_rs2_21_) );
	NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__22_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5681_) );
	MUX2X1 MUX2X1_108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__22_), .B(csr_gpr_iu_gpr_29__22_), .S(biu_ins_20_bF_buf5), .Y(_5682_) );
	OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(_4911__bF_buf4), .C(_5681_), .Y(_5683_) );
	NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf1), .B(_5683_), .Y(_5684_) );
	NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__22_), .B(_4881__bF_buf1), .Y(_5685_) );
	OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_4363_), .B(_4899__bF_buf14), .C(_5685_), .Y(_5686_) );
	OAI22X1 OAI22X1_540 ( .gnd(gnd), .vdd(vdd), .A(_4367_), .B(_4896__bF_buf8), .C(_4366_), .D(_4897__bF_buf14), .Y(_5687_) );
	OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_5687_), .B(_5686_), .C(_4903__bF_buf8), .Y(_5688_) );
	NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf3), .B(_5688_), .C(_5684_), .Y(_5689_) );
	NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__22_), .B(_4881__bF_buf0), .Y(_5690_) );
	OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_2841_), .B(_4897__bF_buf13), .C(_5690_), .Y(_5691_) );
	OAI22X1 OAI22X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .B(_4896__bF_buf7), .C(_2776_), .D(_4899__bF_buf13), .Y(_5692_) );
	OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_5692_), .B(_5691_), .C(_4895__bF_buf0), .Y(_5693_) );
	NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__22_), .B(_4881__bF_buf11), .Y(_5694_) );
	OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_4375_), .B(_4897__bF_buf12), .C(_5694_), .Y(_5695_) );
	OAI22X1 OAI22X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .B(_4896__bF_buf6), .C(_4376_), .D(_4899__bF_buf12), .Y(_5696_) );
	OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_5696_), .B(_5695_), .C(_4903__bF_buf7), .Y(_5697_) );
	NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_5693_), .B(_5697_), .C(_4893__bF_buf2), .Y(_5698_) );
	NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5698_), .C(_5689_), .Y(_5699_) );
	OAI22X1 OAI22X1_543 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .B(_4896__bF_buf5), .C(_4346_), .D(_4897__bF_buf11), .Y(_5700_) );
	NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__22_), .B(_4881__bF_buf10), .Y(_5701_) );
	OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_4899__bF_buf11), .C(_5701_), .Y(_5702_) );
	OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_5700_), .B(_5702_), .C(_4895__bF_buf10), .Y(_5703_) );
	NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__22_), .B(_4881__bF_buf9), .Y(_5704_) );
	OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4899__bF_buf10), .C(_5704_), .Y(_5705_) );
	OAI22X1 OAI22X1_544 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_4896__bF_buf4), .C(_4353_), .D(_4897__bF_buf10), .Y(_5706_) );
	OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_5706_), .B(_5705_), .C(_4903__bF_buf6), .Y(_5707_) );
	AOI22X1 AOI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5703_), .D(_5707_), .Y(_5708_) );
	OAI22X1 OAI22X1_545 ( .gnd(gnd), .vdd(vdd), .A(_4328_), .B(_4896__bF_buf3), .C(_4331_), .D(_4897__bF_buf9), .Y(_5709_) );
	NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__22_), .B(_4881__bF_buf8), .Y(_5710_) );
	OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_4899__bF_buf9), .C(_5710_), .Y(_5711_) );
	OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_5709_), .B(_5711_), .C(_4895__bF_buf9), .Y(_5712_) );
	OAI22X1 OAI22X1_546 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_4896__bF_buf2), .C(_4338_), .D(_4897__bF_buf8), .Y(_5713_) );
	NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__22_), .B(_4881__bF_buf7), .Y(_5714_) );
	OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_4339_), .B(_4899__bF_buf8), .C(_5714_), .Y(_5715_) );
	OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_5713_), .B(_5715_), .C(_4903__bF_buf5), .Y(_5716_) );
	AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_5712_), .B(_5716_), .C(_4893__bF_buf1), .Y(_5717_) );
	OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_5708_), .B(_5717_), .C(_4931__bF_buf2), .Y(_5718_) );
	AOI22X1 AOI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5699_), .D(_5718_), .Y(csr_gpr_iu_rs2_22_) );
	OAI22X1 OAI22X1_547 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(_4896__bF_buf1), .C(_4383_), .D(_4891__bF_buf4), .Y(_5719_) );
	OAI22X1 OAI22X1_548 ( .gnd(gnd), .vdd(vdd), .A(_4386_), .B(_4897__bF_buf7), .C(_4387_), .D(_4899__bF_buf7), .Y(_5720_) );
	OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_5719_), .B(_5720_), .C(_4895__bF_buf8), .Y(_5721_) );
	OAI22X1 OAI22X1_549 ( .gnd(gnd), .vdd(vdd), .A(_4391_), .B(_4896__bF_buf0), .C(_4390_), .D(_4891__bF_buf3), .Y(_5722_) );
	OAI22X1 OAI22X1_550 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_4897__bF_buf6), .C(_4394_), .D(_4899__bF_buf6), .Y(_5723_) );
	OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_5722_), .B(_5723_), .C(_4903__bF_buf4), .Y(_5724_) );
	AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_5724_), .B(_5721_), .C(_4893__bF_buf0), .Y(_5725_) );
	OAI22X1 OAI22X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_4897__bF_buf5), .C(_4398_), .D(_4899__bF_buf5), .Y(_5726_) );
	OAI22X1 OAI22X1_552 ( .gnd(gnd), .vdd(vdd), .A(_4399_), .B(_4896__bF_buf13), .C(_4402_), .D(_4891__bF_buf2), .Y(_5727_) );
	OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_5727_), .B(_5726_), .C(_4895__bF_buf7), .Y(_5728_) );
	OAI22X1 OAI22X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4408_), .B(_4897__bF_buf4), .C(_4405_), .D(_4899__bF_buf4), .Y(_5729_) );
	OAI22X1 OAI22X1_554 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_4896__bF_buf12), .C(_4409_), .D(_4891__bF_buf1), .Y(_5730_) );
	OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_5730_), .B(_5729_), .C(_4903__bF_buf3), .Y(_5731_) );
	AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_5731_), .B(_5728_), .C(_4910__bF_buf2), .Y(_5732_) );
	OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_5732_), .C(_4931__bF_buf1), .Y(_5733_) );
	OAI22X1 OAI22X1_555 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_4897__bF_buf3), .C(_4415_), .D(_4899__bF_buf3), .Y(_5734_) );
	NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__23_), .B(biu_ins_20_bF_buf4), .Y(_5735_) );
	OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(_4417_), .C(_5735_), .Y(_5736_) );
	AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf3), .B(_5736_), .C(_5734_), .Y(_5737_) );
	OAI22X1 OAI22X1_556 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .B(_4897__bF_buf2), .C(_4422_), .D(_4899__bF_buf2), .Y(_5738_) );
	AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__23_), .B(_4911__bF_buf2), .C(_5738_), .Y(_5739_) );
	MUX2X1 MUX2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(_5737_), .S(_4895__bF_buf6), .Y(_5740_) );
	NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__23_), .B(_4881__bF_buf6), .Y(_5741_) );
	OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_2843_), .B(_4897__bF_buf1), .C(_5741_), .Y(_5742_) );
	OAI22X1 OAI22X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_4896__bF_buf11), .C(_2778_), .D(_4899__bF_buf1), .Y(_5743_) );
	OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_5743_), .B(_5742_), .C(_4895__bF_buf5), .Y(_5744_) );
	OAI22X1 OAI22X1_558 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_4897__bF_buf0), .C(_4431_), .D(_4899__bF_buf0), .Y(_5745_) );
	OAI22X1 OAI22X1_559 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_4896__bF_buf10), .C(_4433_), .D(_4891__bF_buf0), .Y(_5746_) );
	OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_5746_), .B(_5745_), .C(_4903__bF_buf2), .Y(_5747_) );
	AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_5744_), .B(_5747_), .C(_4910__bF_buf1), .Y(_5748_) );
	AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_5740_), .B(_4910__bF_buf0), .C(_5748_), .Y(_5749_) );
	OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf3), .B(_5749_), .C(_5733_), .Y(csr_gpr_iu_rs2_23_) );
	NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__24_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5750_) );
	MUX2X1 MUX2X1_110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__24_), .B(csr_gpr_iu_gpr_29__24_), .S(biu_ins_20_bF_buf2), .Y(_5751_) );
	OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_5751_), .B(_4911__bF_buf1), .C(_5750_), .Y(_5752_) );
	NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf4), .B(_5752_), .Y(_5753_) );
	NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__24_), .B(_4881__bF_buf5), .Y(_5754_) );
	OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4899__bF_buf14), .C(_5754_), .Y(_5755_) );
	OAI22X1 OAI22X1_560 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_4896__bF_buf9), .C(_4445_), .D(_4897__bF_buf14), .Y(_5756_) );
	OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_5756_), .B(_5755_), .C(_4903__bF_buf1), .Y(_5757_) );
	NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_5757_), .C(_5753_), .Y(_5758_) );
	OAI22X1 OAI22X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2910_), .B(_4896__bF_buf8), .C(_2845_), .D(_4897__bF_buf13), .Y(_5759_) );
	NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__24_), .B(_4881__bF_buf4), .Y(_5760_) );
	OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_4899__bF_buf13), .C(_5760_), .Y(_5761_) );
	OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_5761_), .C(_4895__bF_buf3), .Y(_5762_) );
	OAI22X1 OAI22X1_562 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_4896__bF_buf7), .C(_4454_), .D(_4897__bF_buf12), .Y(_5763_) );
	NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__24_), .B(_4881__bF_buf3), .Y(_5764_) );
	OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_4899__bF_buf12), .C(_5764_), .Y(_5765_) );
	OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_5763_), .B(_5765_), .C(_4903__bF_buf0), .Y(_5766_) );
	NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_5762_), .B(_5766_), .C(_4893__bF_buf5), .Y(_5767_) );
	NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5767_), .C(_5758_), .Y(_5768_) );
	NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__24_), .B(_4881__bF_buf2), .Y(_5769_) );
	OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_4462_), .B(_4897__bF_buf11), .C(_5769_), .Y(_5770_) );
	OAI22X1 OAI22X1_563 ( .gnd(gnd), .vdd(vdd), .A(_4466_), .B(_4896__bF_buf6), .C(_4465_), .D(_4899__bF_buf11), .Y(_5771_) );
	OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_5771_), .B(_5770_), .C(_4895__bF_buf2), .Y(_5772_) );
	OAI22X1 OAI22X1_564 ( .gnd(gnd), .vdd(vdd), .A(_4473_), .B(_4896__bF_buf5), .C(_4469_), .D(_4899__bF_buf10), .Y(_5773_) );
	NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__24_), .B(_4881__bF_buf1), .Y(_5774_) );
	OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_4472_), .B(_4897__bF_buf10), .C(_5774_), .Y(_5775_) );
	OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_5773_), .B(_5775_), .C(_4903__bF_buf9), .Y(_5776_) );
	AOI22X1 AOI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5772_), .D(_5776_), .Y(_5777_) );
	OAI22X1 OAI22X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_4896__bF_buf4), .C(_4477_), .D(_4897__bF_buf9), .Y(_5778_) );
	NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__24_), .B(_4881__bF_buf0), .Y(_5779_) );
	OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_4899__bF_buf9), .C(_5779_), .Y(_5780_) );
	OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_5778_), .B(_5780_), .C(_4895__bF_buf1), .Y(_5781_) );
	OAI22X1 OAI22X1_566 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_4896__bF_buf3), .C(_4484_), .D(_4897__bF_buf8), .Y(_5782_) );
	NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__24_), .B(_4881__bF_buf11), .Y(_5783_) );
	OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_4899__bF_buf8), .C(_5783_), .Y(_5784_) );
	OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_5782_), .B(_5784_), .C(_4903__bF_buf8), .Y(_5785_) );
	AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(_5785_), .C(_4893__bF_buf4), .Y(_5786_) );
	OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_5777_), .B(_5786_), .C(_4931__bF_buf0), .Y(_5787_) );
	AOI22X1 AOI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5768_), .D(_5787_), .Y(csr_gpr_iu_rs2_24_) );
	NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__25_), .B(_4899__bF_buf7), .C(_4897__bF_buf7), .Y(_5788_) );
	MUX2X1 MUX2X1_111 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__25_), .B(csr_gpr_iu_gpr_29__25_), .S(biu_ins_20_bF_buf1), .Y(_5789_) );
	OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_5789_), .B(_4911__bF_buf0), .C(_5788_), .Y(_5790_) );
	NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf0), .B(_5790_), .Y(_5791_) );
	NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__25_), .B(_4881__bF_buf10), .Y(_5792_) );
	OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_4497_), .B(_4899__bF_buf6), .C(_5792_), .Y(_5793_) );
	OAI22X1 OAI22X1_567 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_4896__bF_buf2), .C(_4500_), .D(_4897__bF_buf6), .Y(_5794_) );
	OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_5794_), .B(_5793_), .C(_4903__bF_buf7), .Y(_5795_) );
	NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf6), .B(_5795_), .C(_5791_), .Y(_5796_) );
	NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__25_), .B(_4881__bF_buf9), .Y(_5797_) );
	OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_4897__bF_buf5), .C(_5797_), .Y(_5798_) );
	OAI22X1 OAI22X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_4896__bF_buf1), .C(_2782_), .D(_4899__bF_buf5), .Y(_5799_) );
	OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_5799_), .B(_5798_), .C(_4895__bF_buf10), .Y(_5800_) );
	NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__25_), .B(_4881__bF_buf8), .Y(_5801_) );
	OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_4509_), .B(_4897__bF_buf4), .C(_5801_), .Y(_5802_) );
	OAI22X1 OAI22X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3045_), .B(_4896__bF_buf0), .C(_4512_), .D(_4899__bF_buf4), .Y(_5803_) );
	OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_5803_), .B(_5802_), .C(_4903__bF_buf6), .Y(_5804_) );
	NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_5800_), .B(_5804_), .C(_4893__bF_buf3), .Y(_5805_) );
	NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5805_), .C(_5796_), .Y(_5806_) );
	OAI22X1 OAI22X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4521_), .B(_4896__bF_buf13), .C(_4517_), .D(_4897__bF_buf3), .Y(_5807_) );
	NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__25_), .B(_4881__bF_buf7), .Y(_5808_) );
	OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_4520_), .B(_4899__bF_buf3), .C(_5808_), .Y(_5809_) );
	OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_5807_), .B(_5809_), .C(_4895__bF_buf9), .Y(_5810_) );
	OAI22X1 OAI22X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4528_), .B(_4896__bF_buf12), .C(_4524_), .D(_4899__bF_buf2), .Y(_5811_) );
	NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__25_), .B(_4881__bF_buf6), .Y(_5812_) );
	OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_4527_), .B(_4897__bF_buf2), .C(_5812_), .Y(_5813_) );
	OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_5813_), .C(_4903__bF_buf5), .Y(_5814_) );
	AOI22X1 AOI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5810_), .D(_5814_), .Y(_5815_) );
	NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__25_), .B(_4881__bF_buf5), .Y(_5816_) );
	OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_4532_), .B(_4897__bF_buf1), .C(_5816_), .Y(_5817_) );
	OAI22X1 OAI22X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_4896__bF_buf11), .C(_4535_), .D(_4899__bF_buf1), .Y(_5818_) );
	OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .B(_5817_), .C(_4895__bF_buf8), .Y(_5819_) );
	NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__25_), .B(_4881__bF_buf4), .Y(_5820_) );
	OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_4897__bF_buf0), .C(_5820_), .Y(_5821_) );
	OAI22X1 OAI22X1_573 ( .gnd(gnd), .vdd(vdd), .A(_4543_), .B(_4896__bF_buf10), .C(_4542_), .D(_4899__bF_buf0), .Y(_5822_) );
	OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_5822_), .B(_5821_), .C(_4903__bF_buf4), .Y(_5823_) );
	AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5823_), .C(_4893__bF_buf2), .Y(_5824_) );
	OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_5815_), .B(_5824_), .C(_4931__bF_buf4), .Y(_5825_) );
	AOI22X1 AOI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5806_), .D(_5825_), .Y(csr_gpr_iu_rs2_25_) );
	OAI22X1 OAI22X1_574 ( .gnd(gnd), .vdd(vdd), .A(_4549_), .B(_4896__bF_buf9), .C(_4548_), .D(_4891__bF_buf7), .Y(_5826_) );
	OAI22X1 OAI22X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_4897__bF_buf15), .C(_4552_), .D(_4899__bF_buf15), .Y(_5827_) );
	OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_5826_), .B(_5827_), .C(_4895__bF_buf7), .Y(_5828_) );
	OAI22X1 OAI22X1_576 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_4896__bF_buf8), .C(_4555_), .D(_4891__bF_buf6), .Y(_5829_) );
	OAI22X1 OAI22X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4558_), .B(_4897__bF_buf14), .C(_4559_), .D(_4899__bF_buf14), .Y(_5830_) );
	OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_5829_), .B(_5830_), .C(_4903__bF_buf3), .Y(_5831_) );
	AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_5831_), .B(_5828_), .C(_4893__bF_buf1), .Y(_5832_) );
	OAI22X1 OAI22X1_578 ( .gnd(gnd), .vdd(vdd), .A(_4566_), .B(_4897__bF_buf13), .C(_4563_), .D(_4899__bF_buf13), .Y(_5833_) );
	OAI22X1 OAI22X1_579 ( .gnd(gnd), .vdd(vdd), .A(_4564_), .B(_4896__bF_buf7), .C(_4567_), .D(_4891__bF_buf5), .Y(_5834_) );
	OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_5834_), .B(_5833_), .C(_4895__bF_buf6), .Y(_5835_) );
	OAI22X1 OAI22X1_580 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_4897__bF_buf12), .C(_4570_), .D(_4899__bF_buf12), .Y(_5836_) );
	OAI22X1 OAI22X1_581 ( .gnd(gnd), .vdd(vdd), .A(_4571_), .B(_4896__bF_buf6), .C(_4574_), .D(_4891__bF_buf4), .Y(_5837_) );
	OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_5837_), .B(_5836_), .C(_4903__bF_buf2), .Y(_5838_) );
	AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_5838_), .B(_5835_), .C(_4910__bF_buf5), .Y(_5839_) );
	OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_5832_), .B(_5839_), .C(_4931__bF_buf3), .Y(_5840_) );
	OAI22X1 OAI22X1_582 ( .gnd(gnd), .vdd(vdd), .A(_4579_), .B(_4897__bF_buf11), .C(_4580_), .D(_4899__bF_buf11), .Y(_5841_) );
	NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__26_), .B(biu_ins_20_bF_buf0), .Y(_5842_) );
	OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf6), .B(_4582_), .C(_5842_), .Y(_5843_) );
	AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf5), .B(_5843_), .C(_5841_), .Y(_5844_) );
	OAI22X1 OAI22X1_583 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4897__bF_buf10), .C(_4587_), .D(_4899__bF_buf10), .Y(_5845_) );
	AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__26_), .B(_4911__bF_buf4), .C(_5845_), .Y(_5846_) );
	MUX2X1 MUX2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_5846_), .B(_5844_), .S(_4895__bF_buf5), .Y(_5847_) );
	NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__26_), .B(_4881__bF_buf3), .Y(_5848_) );
	OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_4897__bF_buf9), .C(_5848_), .Y(_5849_) );
	OAI22X1 OAI22X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_4896__bF_buf5), .C(_2784_), .D(_4899__bF_buf9), .Y(_5850_) );
	OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_5850_), .B(_5849_), .C(_4895__bF_buf4), .Y(_5851_) );
	OAI22X1 OAI22X1_585 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_4897__bF_buf8), .C(_4596_), .D(_4899__bF_buf8), .Y(_5852_) );
	OAI22X1 OAI22X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_4896__bF_buf4), .C(_4598_), .D(_4891__bF_buf3), .Y(_5853_) );
	OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_5853_), .B(_5852_), .C(_4903__bF_buf1), .Y(_5854_) );
	AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_5851_), .B(_5854_), .C(_4910__bF_buf4), .Y(_5855_) );
	AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_5847_), .B(_4910__bF_buf3), .C(_5855_), .Y(_5856_) );
	OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf2), .B(_5856_), .C(_5840_), .Y(csr_gpr_iu_rs2_26_) );
	OAI22X1 OAI22X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .B(_4896__bF_buf3), .C(_4603_), .D(_4891__bF_buf2), .Y(_5857_) );
	OAI22X1 OAI22X1_588 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_4897__bF_buf7), .C(_4607_), .D(_4899__bF_buf7), .Y(_5858_) );
	OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_5857_), .B(_5858_), .C(_4895__bF_buf3), .Y(_5859_) );
	OAI22X1 OAI22X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4896__bF_buf2), .C(_4610_), .D(_4891__bF_buf1), .Y(_5860_) );
	OAI22X1 OAI22X1_590 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_4897__bF_buf6), .C(_4614_), .D(_4899__bF_buf6), .Y(_5861_) );
	OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_5860_), .B(_5861_), .C(_4903__bF_buf0), .Y(_5862_) );
	AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_5862_), .B(_5859_), .C(_4893__bF_buf0), .Y(_5863_) );
	NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__27_), .B(_4881__bF_buf2), .Y(_5864_) );
	OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .B(_4899__bF_buf5), .C(_5864_), .Y(_5865_) );
	OAI22X1 OAI22X1_591 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_4896__bF_buf1), .C(_4618_), .D(_4897__bF_buf5), .Y(_5866_) );
	OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_5866_), .B(_5865_), .C(_4895__bF_buf2), .Y(_5867_) );
	NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__27_), .B(_4881__bF_buf1), .Y(_5868_) );
	OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_4626_), .B(_4899__bF_buf4), .C(_5868_), .Y(_5869_) );
	OAI22X1 OAI22X1_592 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_4896__bF_buf0), .C(_4625_), .D(_4897__bF_buf4), .Y(_5870_) );
	OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_5870_), .B(_5869_), .C(_4903__bF_buf9), .Y(_5871_) );
	AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_5867_), .B(_5871_), .C(_4910__bF_buf2), .Y(_5872_) );
	OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_5863_), .B(_5872_), .C(_4931__bF_buf2), .Y(_5873_) );
	OAI22X1 OAI22X1_593 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_4897__bF_buf3), .C(_4635_), .D(_4899__bF_buf3), .Y(_5874_) );
	NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__27_), .B(biu_ins_20_bF_buf5), .Y(_5875_) );
	OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf4), .B(_4637_), .C(_5875_), .Y(_5876_) );
	AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf3), .B(_5876_), .C(_5874_), .Y(_5877_) );
	OAI22X1 OAI22X1_594 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .B(_4897__bF_buf2), .C(_4642_), .D(_4899__bF_buf2), .Y(_5878_) );
	AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__27_), .B(_4911__bF_buf2), .C(_5878_), .Y(_5879_) );
	MUX2X1 MUX2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_5879_), .B(_5877_), .S(_4895__bF_buf1), .Y(_5880_) );
	NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__27_), .B(_4881__bF_buf0), .Y(_5881_) );
	OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_2851_), .B(_4897__bF_buf1), .C(_5881_), .Y(_5882_) );
	OAI22X1 OAI22X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .B(_4896__bF_buf13), .C(_2786_), .D(_4899__bF_buf1), .Y(_5883_) );
	OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_5882_), .C(_4895__bF_buf0), .Y(_5884_) );
	OAI22X1 OAI22X1_596 ( .gnd(gnd), .vdd(vdd), .A(_4650_), .B(_4897__bF_buf0), .C(_4651_), .D(_4899__bF_buf0), .Y(_5885_) );
	OAI22X1 OAI22X1_597 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_4896__bF_buf12), .C(_4653_), .D(_4891__bF_buf0), .Y(_5886_) );
	OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .B(_5885_), .C(_4903__bF_buf8), .Y(_5887_) );
	AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_5887_), .C(_4910__bF_buf1), .Y(_5888_) );
	AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_5880_), .B(_4910__bF_buf0), .C(_5888_), .Y(_5889_) );
	OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf1), .B(_5889_), .C(_5873_), .Y(csr_gpr_iu_rs2_27_) );
	NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__28_), .B(_4899__bF_buf15), .C(_4897__bF_buf15), .Y(_5890_) );
	MUX2X1 MUX2X1_114 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__28_), .B(csr_gpr_iu_gpr_29__28_), .S(biu_ins_20_bF_buf3), .Y(_5891_) );
	OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_5891_), .B(_4911__bF_buf1), .C(_5890_), .Y(_5892_) );
	NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_4895__bF_buf10), .B(_5892_), .Y(_5893_) );
	NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_27__28_), .B(_4881__bF_buf11), .Y(_5894_) );
	OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4899__bF_buf14), .C(_5894_), .Y(_5895_) );
	OAI22X1 OAI22X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4666_), .B(_4896__bF_buf11), .C(_4665_), .D(_4897__bF_buf14), .Y(_5896_) );
	OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_5896_), .B(_5895_), .C(_4903__bF_buf7), .Y(_5897_) );
	NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4910__bF_buf7), .B(_5897_), .C(_5893_), .Y(_5898_) );
	OAI22X1 OAI22X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .B(_4896__bF_buf10), .C(_2853_), .D(_4897__bF_buf13), .Y(_5899_) );
	NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__28_), .B(_4881__bF_buf10), .Y(_5900_) );
	OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_4899__bF_buf13), .C(_5900_), .Y(_5901_) );
	OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_5899_), .B(_5901_), .C(_4895__bF_buf9), .Y(_5902_) );
	OAI22X1 OAI22X1_600 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_4896__bF_buf9), .C(_4674_), .D(_4897__bF_buf12), .Y(_5903_) );
	NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_19__28_), .B(_4881__bF_buf9), .Y(_5904_) );
	OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_4899__bF_buf12), .C(_5904_), .Y(_5905_) );
	OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_5903_), .B(_5905_), .C(_4903__bF_buf6), .Y(_5906_) );
	NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_5902_), .B(_5906_), .C(_4893__bF_buf5), .Y(_5907_) );
	NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5907_), .C(_5898_), .Y(_5908_) );
	OAI22X1 OAI22X1_601 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_4896__bF_buf8), .C(_4682_), .D(_4897__bF_buf11), .Y(_5909_) );
	NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__28_), .B(_4881__bF_buf8), .Y(_5910_) );
	OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_4685_), .B(_4899__bF_buf11), .C(_5910_), .Y(_5911_) );
	OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_5909_), .B(_5911_), .C(_4895__bF_buf8), .Y(_5912_) );
	NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__28_), .B(_4881__bF_buf7), .Y(_5913_) );
	OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_4689_), .B(_4899__bF_buf10), .C(_5913_), .Y(_5914_) );
	OAI22X1 OAI22X1_602 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4896__bF_buf7), .C(_4692_), .D(_4897__bF_buf10), .Y(_5915_) );
	OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .B(_5914_), .C(_4903__bF_buf5), .Y(_5916_) );
	AOI22X1 AOI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4892_), .C(_5912_), .D(_5916_), .Y(_5917_) );
	NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_15__28_), .B(_4881__bF_buf6), .Y(_5918_) );
	OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_4697_), .B(_4897__bF_buf9), .C(_5918_), .Y(_5919_) );
	OAI22X1 OAI22X1_603 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_4896__bF_buf6), .C(_4700_), .D(_4899__bF_buf9), .Y(_5920_) );
	OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .B(_5919_), .C(_4895__bF_buf7), .Y(_5921_) );
	NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_11__28_), .B(_4881__bF_buf5), .Y(_5922_) );
	OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4897__bF_buf8), .C(_5922_), .Y(_5923_) );
	OAI22X1 OAI22X1_604 ( .gnd(gnd), .vdd(vdd), .A(_4705_), .B(_4896__bF_buf5), .C(_4707_), .D(_4899__bF_buf8), .Y(_5924_) );
	OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_5924_), .B(_5923_), .C(_4903__bF_buf4), .Y(_5925_) );
	AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .B(_5925_), .C(_4893__bF_buf4), .Y(_5926_) );
	OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_5917_), .B(_5926_), .C(_4931__bF_buf1), .Y(_5927_) );
	AOI22X1 AOI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_4883_), .C(_5908_), .D(_5927_), .Y(csr_gpr_iu_rs2_28_) );
	OAI22X1 OAI22X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_4896__bF_buf4), .C(_4753_), .D(_4891__bF_buf7), .Y(_5928_) );
	OAI22X1 OAI22X1_606 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_4897__bF_buf7), .C(_4755_), .D(_4899__bF_buf7), .Y(_5929_) );
	OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_5928_), .B(_5929_), .C(_4895__bF_buf6), .Y(_5930_) );
	OAI22X1 OAI22X1_607 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_4896__bF_buf3), .C(_4760_), .D(_4891__bF_buf6), .Y(_5931_) );
	OAI22X1 OAI22X1_608 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(_4897__bF_buf6), .C(_4762_), .D(_4899__bF_buf6), .Y(_5932_) );
	OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_5931_), .B(_5932_), .C(_4903__bF_buf3), .Y(_5933_) );
	AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_5933_), .B(_5930_), .C(_4893__bF_buf3), .Y(_5934_) );
	OAI22X1 OAI22X1_609 ( .gnd(gnd), .vdd(vdd), .A(_4737_), .B(_4897__bF_buf5), .C(_4740_), .D(_4899__bF_buf5), .Y(_5935_) );
	OAI22X1 OAI22X1_610 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_4896__bF_buf2), .C(_4741_), .D(_4891__bF_buf5), .Y(_5936_) );
	OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_5936_), .B(_5935_), .C(_4895__bF_buf5), .Y(_5937_) );
	OAI22X1 OAI22X1_611 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(_4897__bF_buf4), .C(_4744_), .D(_4899__bF_buf4), .Y(_5938_) );
	OAI22X1 OAI22X1_612 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_4896__bF_buf1), .C(_4748_), .D(_4891__bF_buf4), .Y(_5939_) );
	OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_5939_), .B(_5938_), .C(_4903__bF_buf2), .Y(_5940_) );
	AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_5940_), .B(_5937_), .C(_4910__bF_buf6), .Y(_5941_) );
	OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_5934_), .B(_5941_), .C(_4931__bF_buf0), .Y(_5942_) );
	INVX1 INVX1_1111 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_29__29_), .Y(_5943_) );
	INVX1 INVX1_1112 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_28__29_), .Y(_5944_) );
	OAI22X1 OAI22X1_613 ( .gnd(gnd), .vdd(vdd), .A(_5943_), .B(_4897__bF_buf3), .C(_5944_), .D(_4899__bF_buf3), .Y(_5945_) );
	AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__29_), .B(_4911__bF_buf0), .C(_5945_), .Y(_5946_) );
	OAI22X1 OAI22X1_614 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_4899__bF_buf2), .C(_4717_), .D(_4891__bF_buf3), .Y(_5947_) );
	OAI22X1 OAI22X1_615 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_4896__bF_buf0), .C(_4720_), .D(_4897__bF_buf2), .Y(_5948_) );
	OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_5947_), .B(_5948_), .C(_4903__bF_buf1), .Y(_5949_) );
	OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_4903__bF_buf0), .B(_5946_), .C(_5949_), .Y(_5950_) );
	NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__29_), .B(_4881__bF_buf4), .Y(_5951_) );
	OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_4897__bF_buf1), .C(_5951_), .Y(_5952_) );
	OAI22X1 OAI22X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_4896__bF_buf13), .C(_2790_), .D(_4899__bF_buf1), .Y(_5953_) );
	OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .B(_5952_), .C(_4895__bF_buf4), .Y(_5954_) );
	OAI22X1 OAI22X1_617 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_4897__bF_buf0), .C(_4732_), .D(_4899__bF_buf0), .Y(_5955_) );
	OAI22X1 OAI22X1_618 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_4896__bF_buf12), .C(_4731_), .D(_4891__bF_buf2), .Y(_5956_) );
	OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_5956_), .B(_5955_), .C(_4903__bF_buf9), .Y(_5957_) );
	AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_5954_), .B(_5957_), .C(_4910__bF_buf5), .Y(_5958_) );
	AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_5950_), .B(_4910__bF_buf4), .C(_5958_), .Y(_5959_) );
	OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf0), .B(_5959_), .C(_5942_), .Y(csr_gpr_iu_rs2_29_) );
	OAI22X1 OAI22X1_619 ( .gnd(gnd), .vdd(vdd), .A(_4769_), .B(_4896__bF_buf11), .C(_4768_), .D(_4891__bF_buf1), .Y(_5960_) );
	OAI22X1 OAI22X1_620 ( .gnd(gnd), .vdd(vdd), .A(_4771_), .B(_4897__bF_buf15), .C(_4772_), .D(_4899__bF_buf15), .Y(_5961_) );
	OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_5960_), .B(_5961_), .C(_4895__bF_buf3), .Y(_5962_) );
	OAI22X1 OAI22X1_621 ( .gnd(gnd), .vdd(vdd), .A(_4776_), .B(_4896__bF_buf10), .C(_4775_), .D(_4891__bF_buf0), .Y(_5963_) );
	OAI22X1 OAI22X1_622 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_4897__bF_buf14), .C(_4779_), .D(_4899__bF_buf14), .Y(_5964_) );
	OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_5963_), .B(_5964_), .C(_4903__bF_buf8), .Y(_5965_) );
	AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_5965_), .B(_5962_), .C(_4893__bF_buf2), .Y(_5966_) );
	NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_7__30_), .B(_4881__bF_buf3), .Y(_5967_) );
	OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4899__bF_buf13), .C(_5967_), .Y(_5968_) );
	OAI22X1 OAI22X1_623 ( .gnd(gnd), .vdd(vdd), .A(_4784_), .B(_4896__bF_buf9), .C(_4786_), .D(_4897__bF_buf13), .Y(_5969_) );
	OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_5969_), .B(_5968_), .C(_4895__bF_buf2), .Y(_5970_) );
	NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_3__30_), .B(_4881__bF_buf2), .Y(_5971_) );
	OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4899__bF_buf12), .C(_5971_), .Y(_5972_) );
	OAI22X1 OAI22X1_624 ( .gnd(gnd), .vdd(vdd), .A(_4791_), .B(_4896__bF_buf8), .C(_4793_), .D(_4897__bF_buf12), .Y(_5973_) );
	OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_5973_), .B(_5972_), .C(_4903__bF_buf7), .Y(_5974_) );
	AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .B(_5974_), .C(_4910__bF_buf3), .Y(_5975_) );
	OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_5966_), .B(_5975_), .C(_4931__bF_buf4), .Y(_5976_) );
	OAI22X1 OAI22X1_625 ( .gnd(gnd), .vdd(vdd), .A(_4799_), .B(_4897__bF_buf11), .C(_4800_), .D(_4899__bF_buf11), .Y(_5977_) );
	NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__30_), .B(biu_ins_20_bF_buf2), .Y(_5978_) );
	OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf1), .B(_4802_), .C(_5978_), .Y(_5979_) );
	AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf5), .B(_5979_), .C(_5977_), .Y(_5980_) );
	OAI22X1 OAI22X1_626 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(_4897__bF_buf10), .C(_4807_), .D(_4899__bF_buf10), .Y(_5981_) );
	AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__30_), .B(_4911__bF_buf4), .C(_5981_), .Y(_5982_) );
	MUX2X1 MUX2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_5980_), .S(_4895__bF_buf1), .Y(_5983_) );
	NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__30_), .B(_4881__bF_buf1), .Y(_5984_) );
	OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_4897__bF_buf9), .C(_5984_), .Y(_5985_) );
	OAI22X1 OAI22X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_4896__bF_buf7), .C(_2792_), .D(_4899__bF_buf9), .Y(_5986_) );
	OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_5986_), .B(_5985_), .C(_4895__bF_buf0), .Y(_5987_) );
	OAI22X1 OAI22X1_628 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_4897__bF_buf8), .C(_4816_), .D(_4899__bF_buf8), .Y(_5988_) );
	OAI22X1 OAI22X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_4896__bF_buf6), .C(_4818_), .D(_4891__bF_buf7), .Y(_5989_) );
	OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_5989_), .B(_5988_), .C(_4903__bF_buf6), .Y(_5990_) );
	AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .B(_5990_), .C(_4910__bF_buf2), .Y(_5991_) );
	AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_5983_), .B(_4910__bF_buf1), .C(_5991_), .Y(_5992_) );
	OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf3), .B(_5992_), .C(_5976_), .Y(csr_gpr_iu_rs2_30_) );
	OAI22X1 OAI22X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_4896__bF_buf5), .C(_4823_), .D(_4891__bF_buf6), .Y(_5993_) );
	OAI22X1 OAI22X1_631 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_4897__bF_buf7), .C(_4827_), .D(_4899__bF_buf7), .Y(_5994_) );
	OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_5993_), .B(_5994_), .C(_4895__bF_buf10), .Y(_5995_) );
	OAI22X1 OAI22X1_632 ( .gnd(gnd), .vdd(vdd), .A(_4831_), .B(_4896__bF_buf4), .C(_4830_), .D(_4891__bF_buf5), .Y(_5996_) );
	OAI22X1 OAI22X1_633 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_4897__bF_buf6), .C(_4834_), .D(_4899__bF_buf6), .Y(_5997_) );
	OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(_5997_), .C(_4903__bF_buf5), .Y(_5998_) );
	AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_5998_), .B(_5995_), .C(_4893__bF_buf1), .Y(_5999_) );
	OAI22X1 OAI22X1_634 ( .gnd(gnd), .vdd(vdd), .A(_4841_), .B(_4897__bF_buf5), .C(_4838_), .D(_4899__bF_buf5), .Y(_6000_) );
	OAI22X1 OAI22X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_4896__bF_buf3), .C(_4839_), .D(_4891__bF_buf4), .Y(_6001_) );
	OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_6001_), .B(_6000_), .C(_4895__bF_buf9), .Y(_6002_) );
	OAI22X1 OAI22X1_636 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_4897__bF_buf4), .C(_4845_), .D(_4899__bF_buf4), .Y(_6003_) );
	OAI22X1 OAI22X1_637 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .B(_4896__bF_buf2), .C(_4846_), .D(_4891__bF_buf3), .Y(_6004_) );
	OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_6004_), .B(_6003_), .C(_4903__bF_buf4), .Y(_6005_) );
	AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_6005_), .B(_6002_), .C(_4910__bF_buf0), .Y(_6006_) );
	OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_5999_), .B(_6006_), .C(_4931__bF_buf3), .Y(_6007_) );
	OAI22X1 OAI22X1_638 ( .gnd(gnd), .vdd(vdd), .A(_4854_), .B(_4897__bF_buf3), .C(_4855_), .D(_4899__bF_buf3), .Y(_6008_) );
	NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_26__31_), .B(biu_ins_20_bF_buf0), .Y(_6009_) );
	OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf6), .B(_4857_), .C(_6009_), .Y(_6010_) );
	AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_4911__bF_buf3), .B(_6010_), .C(_6008_), .Y(_6011_) );
	OAI22X1 OAI22X1_639 ( .gnd(gnd), .vdd(vdd), .A(_4861_), .B(_4897__bF_buf2), .C(_4862_), .D(_4899__bF_buf2), .Y(_6012_) );
	AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_30__31_), .B(_4911__bF_buf2), .C(_6012_), .Y(_6013_) );
	MUX2X1 MUX2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_6013_), .B(_6011_), .S(_4895__bF_buf8), .Y(_6014_) );
	OAI22X1 OAI22X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_4896__bF_buf1), .C(_2859_), .D(_4897__bF_buf1), .Y(_6015_) );
	NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_gpr_23__31_), .B(_4881__bF_buf0), .Y(_6016_) );
	OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .B(_4899__bF_buf1), .C(_6016_), .Y(_6017_) );
	OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_6015_), .B(_6017_), .C(_4895__bF_buf7), .Y(_6018_) );
	OAI22X1 OAI22X1_641 ( .gnd(gnd), .vdd(vdd), .A(_4870_), .B(_4897__bF_buf0), .C(_4871_), .D(_4899__bF_buf0), .Y(_6019_) );
	OAI22X1 OAI22X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .B(_4896__bF_buf0), .C(_4873_), .D(_4891__bF_buf2), .Y(_6020_) );
	OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_6020_), .B(_6019_), .C(_4903__bF_buf3), .Y(_6021_) );
	AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_6018_), .B(_6021_), .C(_4910__bF_buf7), .Y(_6022_) );
	AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_4910__bF_buf6), .C(_6022_), .Y(_6023_) );
	OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_4886__bF_buf2), .B(_6023_), .C(_6007_), .Y(csr_gpr_iu_rs2_31_) );
	AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_2476_), .B(_2486_), .Y(_6024_) );
	NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2588__bF_buf5), .C(_6024_), .Y(_6025_) );
	NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2482_), .C(_2476_), .Y(_6026_) );
	OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2590__bF_buf11), .C(csr_gpr_iu_gpr_14__0_), .Y(_6027_) );
	OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf0), .B(_6025__bF_buf4), .C(_6027_), .Y(_1756_) );
	OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2590__bF_buf10), .C(csr_gpr_iu_gpr_14__1_), .Y(_6028_) );
	OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf0), .B(_6025__bF_buf3), .C(_6028_), .Y(_1757_) );
	OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2590__bF_buf9), .C(csr_gpr_iu_gpr_14__2_), .Y(_6029_) );
	OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf0), .B(_6025__bF_buf2), .C(_6029_), .Y(_1758_) );
	OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2590__bF_buf8), .C(csr_gpr_iu_gpr_14__3_), .Y(_6030_) );
	OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf0), .B(_6025__bF_buf1), .C(_6030_), .Y(_1759_) );
	OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2590__bF_buf7), .C(csr_gpr_iu_gpr_14__4_), .Y(_6031_) );
	OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf0), .B(_6025__bF_buf0), .C(_6031_), .Y(_1760_) );
	OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_14__5_), .Y(_6032_) );
	OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf0), .B(_6025__bF_buf4), .C(_6032_), .Y(_1761_) );
	OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2590__bF_buf5), .C(csr_gpr_iu_gpr_14__6_), .Y(_6033_) );
	OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf0), .B(_6025__bF_buf3), .C(_6033_), .Y(_1762_) );
	OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2590__bF_buf4), .C(csr_gpr_iu_gpr_14__7_), .Y(_6034_) );
	OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf0), .B(_6025__bF_buf2), .C(_6034_), .Y(_1763_) );
	OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2590__bF_buf3), .C(csr_gpr_iu_gpr_14__8_), .Y(_6035_) );
	OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf0), .B(_6025__bF_buf1), .C(_6035_), .Y(_1764_) );
	OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2590__bF_buf2), .C(csr_gpr_iu_gpr_14__9_), .Y(_6036_) );
	OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf0), .B(_6025__bF_buf0), .C(_6036_), .Y(_1765_) );
	OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2590__bF_buf1), .C(csr_gpr_iu_gpr_14__10_), .Y(_6037_) );
	OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf0), .B(_6025__bF_buf4), .C(_6037_), .Y(_1766_) );
	OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2590__bF_buf0), .C(csr_gpr_iu_gpr_14__11_), .Y(_6038_) );
	OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf0), .B(_6025__bF_buf3), .C(_6038_), .Y(_1767_) );
	OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2590__bF_buf12), .C(csr_gpr_iu_gpr_14__12_), .Y(_6039_) );
	OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf0), .B(_6025__bF_buf2), .C(_6039_), .Y(_1768_) );
	OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2590__bF_buf11), .C(csr_gpr_iu_gpr_14__13_), .Y(_6040_) );
	OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf0), .B(_6025__bF_buf1), .C(_6040_), .Y(_1769_) );
	OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2590__bF_buf10), .C(csr_gpr_iu_gpr_14__14_), .Y(_6041_) );
	OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf0), .B(_6025__bF_buf0), .C(_6041_), .Y(_1770_) );
	OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2590__bF_buf9), .C(csr_gpr_iu_gpr_14__15_), .Y(_6042_) );
	OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf0), .B(_6025__bF_buf4), .C(_6042_), .Y(_1771_) );
	OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2590__bF_buf8), .C(csr_gpr_iu_gpr_14__16_), .Y(_6043_) );
	OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf0), .B(_6025__bF_buf3), .C(_6043_), .Y(_1772_) );
	OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2590__bF_buf7), .C(csr_gpr_iu_gpr_14__17_), .Y(_6044_) );
	OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf0), .B(_6025__bF_buf2), .C(_6044_), .Y(_1773_) );
	OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_14__18_), .Y(_6045_) );
	OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf0), .B(_6025__bF_buf1), .C(_6045_), .Y(_1774_) );
	OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2590__bF_buf5), .C(csr_gpr_iu_gpr_14__19_), .Y(_6046_) );
	OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf0), .B(_6025__bF_buf0), .C(_6046_), .Y(_1775_) );
	OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2590__bF_buf4), .C(csr_gpr_iu_gpr_14__20_), .Y(_6047_) );
	OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf0), .B(_6025__bF_buf4), .C(_6047_), .Y(_1776_) );
	OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2590__bF_buf3), .C(csr_gpr_iu_gpr_14__21_), .Y(_6048_) );
	OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf0), .B(_6025__bF_buf3), .C(_6048_), .Y(_1777_) );
	OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2590__bF_buf2), .C(csr_gpr_iu_gpr_14__22_), .Y(_6049_) );
	OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf0), .B(_6025__bF_buf2), .C(_6049_), .Y(_1778_) );
	OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2590__bF_buf1), .C(csr_gpr_iu_gpr_14__23_), .Y(_6050_) );
	OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf0), .B(_6025__bF_buf1), .C(_6050_), .Y(_1779_) );
	OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2590__bF_buf0), .C(csr_gpr_iu_gpr_14__24_), .Y(_6051_) );
	OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf0), .B(_6025__bF_buf0), .C(_6051_), .Y(_1780_) );
	OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2590__bF_buf12), .C(csr_gpr_iu_gpr_14__25_), .Y(_6052_) );
	OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf0), .B(_6025__bF_buf4), .C(_6052_), .Y(_1781_) );
	OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2590__bF_buf11), .C(csr_gpr_iu_gpr_14__26_), .Y(_6053_) );
	OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf0), .B(_6025__bF_buf3), .C(_6053_), .Y(_1782_) );
	OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2590__bF_buf10), .C(csr_gpr_iu_gpr_14__27_), .Y(_6054_) );
	OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf0), .B(_6025__bF_buf2), .C(_6054_), .Y(_1783_) );
	OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2590__bF_buf9), .C(csr_gpr_iu_gpr_14__28_), .Y(_6055_) );
	OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf0), .B(_6025__bF_buf1), .C(_6055_), .Y(_1784_) );
	OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2590__bF_buf8), .C(csr_gpr_iu_gpr_14__29_), .Y(_6056_) );
	OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf0), .B(_6025__bF_buf0), .C(_6056_), .Y(_1785_) );
	OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2590__bF_buf7), .C(csr_gpr_iu_gpr_14__30_), .Y(_6057_) );
	OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_6025__bF_buf4), .C(_6057_), .Y(_1786_) );
	OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_14__31_), .Y(_6058_) );
	OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf0), .B(_6025__bF_buf3), .C(_6058_), .Y(_1787_) );
	NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf1), .B(_2696__bF_buf12), .Y(_6059_) );
	NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2995__bF_buf2), .C(_2694__bF_buf5), .Y(_6060_) );
	OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_6059__bF_buf4), .C(_6060_), .Y(_1788_) );
	NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2995__bF_buf1), .C(_2694__bF_buf4), .Y(_6061_) );
	OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .B(_6059__bF_buf3), .C(_6061_), .Y(_1789_) );
	NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2995__bF_buf0), .C(_2694__bF_buf3), .Y(_6062_) );
	OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_3276_), .B(_6059__bF_buf2), .C(_6062_), .Y(_1790_) );
	NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2995__bF_buf8), .C(_2694__bF_buf2), .Y(_6063_) );
	OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_6059__bF_buf1), .C(_6063_), .Y(_1791_) );
	NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2995__bF_buf7), .C(_2694__bF_buf1), .Y(_6064_) );
	OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_6059__bF_buf0), .C(_6064_), .Y(_1792_) );
	NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2995__bF_buf6), .C(_2694__bF_buf0), .Y(_6065_) );
	OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_3441_), .B(_6059__bF_buf4), .C(_6065_), .Y(_1793_) );
	NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2995__bF_buf5), .C(_2694__bF_buf7), .Y(_6066_) );
	OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_3496_), .B(_6059__bF_buf3), .C(_6066_), .Y(_1794_) );
	NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2995__bF_buf4), .C(_2694__bF_buf6), .Y(_6067_) );
	OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_3522_), .B(_6059__bF_buf2), .C(_6067_), .Y(_1795_) );
	NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2995__bF_buf3), .C(_2694__bF_buf5), .Y(_6068_) );
	OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .B(_6059__bF_buf1), .C(_6068_), .Y(_1796_) );
	NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2995__bF_buf2), .C(_2694__bF_buf4), .Y(_6069_) );
	OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_6059__bF_buf0), .C(_6069_), .Y(_1797_) );
	NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2995__bF_buf1), .C(_2694__bF_buf3), .Y(_6070_) );
	OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_6059__bF_buf4), .C(_6070_), .Y(_1798_) );
	NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2995__bF_buf0), .C(_2694__bF_buf2), .Y(_6071_) );
	OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_6059__bF_buf3), .C(_6071_), .Y(_1799_) );
	NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2995__bF_buf8), .C(_2694__bF_buf1), .Y(_6072_) );
	OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_6059__bF_buf2), .C(_6072_), .Y(_1800_) );
	NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2995__bF_buf7), .C(_2694__bF_buf0), .Y(_6073_) );
	OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_3881_), .B(_6059__bF_buf1), .C(_6073_), .Y(_1801_) );
	NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2995__bF_buf6), .C(_2694__bF_buf7), .Y(_6074_) );
	OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_6059__bF_buf0), .C(_6074_), .Y(_1802_) );
	NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2995__bF_buf5), .C(_2694__bF_buf6), .Y(_6075_) );
	OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_6059__bF_buf4), .C(_6075_), .Y(_1803_) );
	NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2995__bF_buf4), .C(_2694__bF_buf5), .Y(_6076_) );
	OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_4016_), .B(_6059__bF_buf3), .C(_6076_), .Y(_1804_) );
	NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2995__bF_buf3), .C(_2694__bF_buf4), .Y(_6077_) );
	OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_4072_), .B(_6059__bF_buf2), .C(_6077_), .Y(_1805_) );
	NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2995__bF_buf2), .C(_2694__bF_buf3), .Y(_6078_) );
	OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_4127_), .B(_6059__bF_buf1), .C(_6078_), .Y(_1806_) );
	NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2995__bF_buf1), .C(_2694__bF_buf2), .Y(_6079_) );
	OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_4211_), .B(_6059__bF_buf0), .C(_6079_), .Y(_1807_) );
	NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2995__bF_buf0), .C(_2694__bF_buf1), .Y(_6080_) );
	OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_6059__bF_buf4), .C(_6080_), .Y(_1808_) );
	NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2995__bF_buf8), .C(_2694__bF_buf0), .Y(_6081_) );
	OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .B(_6059__bF_buf3), .C(_6081_), .Y(_1809_) );
	NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2995__bF_buf7), .C(_2694__bF_buf7), .Y(_6082_) );
	OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_4376_), .B(_6059__bF_buf2), .C(_6082_), .Y(_1810_) );
	NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2995__bF_buf6), .C(_2694__bF_buf6), .Y(_6083_) );
	OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_4431_), .B(_6059__bF_buf1), .C(_6083_), .Y(_1811_) );
	NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2995__bF_buf5), .C(_2694__bF_buf5), .Y(_6084_) );
	OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_6059__bF_buf0), .C(_6084_), .Y(_1812_) );
	NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2995__bF_buf4), .C(_2694__bF_buf4), .Y(_6085_) );
	OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_4512_), .B(_6059__bF_buf4), .C(_6085_), .Y(_1813_) );
	NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2995__bF_buf3), .C(_2694__bF_buf3), .Y(_6086_) );
	OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_4596_), .B(_6059__bF_buf3), .C(_6086_), .Y(_1814_) );
	NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2995__bF_buf2), .C(_2694__bF_buf2), .Y(_6087_) );
	OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_6059__bF_buf2), .C(_6087_), .Y(_1815_) );
	NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2995__bF_buf1), .C(_2694__bF_buf1), .Y(_6088_) );
	OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_6059__bF_buf1), .C(_6088_), .Y(_1816_) );
	NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2995__bF_buf0), .C(_2694__bF_buf0), .Y(_6089_) );
	OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(_6059__bF_buf0), .C(_6089_), .Y(_1817_) );
	NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2995__bF_buf8), .C(_2694__bF_buf7), .Y(_6090_) );
	OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .B(_6059__bF_buf4), .C(_6090_), .Y(_1818_) );
	NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2995__bF_buf7), .C(_2694__bF_buf6), .Y(_6091_) );
	OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .B(_6059__bF_buf3), .C(_6091_), .Y(_1819_) );
	OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2625__bF_buf8), .Y(_6092_) );
	OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6026__bF_buf10), .C(csr_gpr_iu_gpr_15__0_), .Y(_6093_) );
	OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf4), .B(_6092__bF_buf4), .C(_6093_), .Y(_1820_) );
	OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6026__bF_buf9), .C(csr_gpr_iu_gpr_15__1_), .Y(_6094_) );
	OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf4), .B(_6092__bF_buf3), .C(_6094_), .Y(_1821_) );
	OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6026__bF_buf8), .C(csr_gpr_iu_gpr_15__2_), .Y(_6095_) );
	OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf4), .B(_6092__bF_buf2), .C(_6095_), .Y(_1822_) );
	OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6026__bF_buf7), .C(csr_gpr_iu_gpr_15__3_), .Y(_6096_) );
	OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf4), .B(_6092__bF_buf1), .C(_6096_), .Y(_1823_) );
	OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6026__bF_buf6), .C(csr_gpr_iu_gpr_15__4_), .Y(_6097_) );
	OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf4), .B(_6092__bF_buf0), .C(_6097_), .Y(_1824_) );
	OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6026__bF_buf5), .C(csr_gpr_iu_gpr_15__5_), .Y(_6098_) );
	OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf4), .B(_6092__bF_buf4), .C(_6098_), .Y(_1825_) );
	OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6026__bF_buf4), .C(csr_gpr_iu_gpr_15__6_), .Y(_6099_) );
	OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf4), .B(_6092__bF_buf3), .C(_6099_), .Y(_1826_) );
	OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6026__bF_buf3), .C(csr_gpr_iu_gpr_15__7_), .Y(_6100_) );
	OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf4), .B(_6092__bF_buf2), .C(_6100_), .Y(_1827_) );
	OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6026__bF_buf2), .C(csr_gpr_iu_gpr_15__8_), .Y(_6101_) );
	OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf4), .B(_6092__bF_buf1), .C(_6101_), .Y(_1828_) );
	OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6026__bF_buf1), .C(csr_gpr_iu_gpr_15__9_), .Y(_6102_) );
	OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf4), .B(_6092__bF_buf0), .C(_6102_), .Y(_1829_) );
	OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6026__bF_buf0), .C(csr_gpr_iu_gpr_15__10_), .Y(_6103_) );
	OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf4), .B(_6092__bF_buf4), .C(_6103_), .Y(_1830_) );
	OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6026__bF_buf10), .C(csr_gpr_iu_gpr_15__11_), .Y(_6104_) );
	OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf4), .B(_6092__bF_buf3), .C(_6104_), .Y(_1831_) );
	OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6026__bF_buf9), .C(csr_gpr_iu_gpr_15__12_), .Y(_6105_) );
	OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf4), .B(_6092__bF_buf2), .C(_6105_), .Y(_1832_) );
	OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6026__bF_buf8), .C(csr_gpr_iu_gpr_15__13_), .Y(_6106_) );
	OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf4), .B(_6092__bF_buf1), .C(_6106_), .Y(_1833_) );
	OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6026__bF_buf7), .C(csr_gpr_iu_gpr_15__14_), .Y(_6107_) );
	OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf4), .B(_6092__bF_buf0), .C(_6107_), .Y(_1834_) );
	OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6026__bF_buf6), .C(csr_gpr_iu_gpr_15__15_), .Y(_6108_) );
	OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf4), .B(_6092__bF_buf4), .C(_6108_), .Y(_1835_) );
	OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6026__bF_buf5), .C(csr_gpr_iu_gpr_15__16_), .Y(_6109_) );
	OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf4), .B(_6092__bF_buf3), .C(_6109_), .Y(_1836_) );
	OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6026__bF_buf4), .C(csr_gpr_iu_gpr_15__17_), .Y(_6110_) );
	OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf4), .B(_6092__bF_buf2), .C(_6110_), .Y(_1837_) );
	OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6026__bF_buf3), .C(csr_gpr_iu_gpr_15__18_), .Y(_6111_) );
	OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf4), .B(_6092__bF_buf1), .C(_6111_), .Y(_1838_) );
	OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6026__bF_buf2), .C(csr_gpr_iu_gpr_15__19_), .Y(_6112_) );
	OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf4), .B(_6092__bF_buf0), .C(_6112_), .Y(_1839_) );
	OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6026__bF_buf1), .C(csr_gpr_iu_gpr_15__20_), .Y(_6113_) );
	OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf4), .B(_6092__bF_buf4), .C(_6113_), .Y(_1840_) );
	OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6026__bF_buf0), .C(csr_gpr_iu_gpr_15__21_), .Y(_6114_) );
	OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf4), .B(_6092__bF_buf3), .C(_6114_), .Y(_1841_) );
	OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6026__bF_buf10), .C(csr_gpr_iu_gpr_15__22_), .Y(_6115_) );
	OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf4), .B(_6092__bF_buf2), .C(_6115_), .Y(_1842_) );
	OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6026__bF_buf9), .C(csr_gpr_iu_gpr_15__23_), .Y(_6116_) );
	OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf4), .B(_6092__bF_buf1), .C(_6116_), .Y(_1843_) );
	OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6026__bF_buf8), .C(csr_gpr_iu_gpr_15__24_), .Y(_6117_) );
	OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf4), .B(_6092__bF_buf0), .C(_6117_), .Y(_1844_) );
	OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6026__bF_buf7), .C(csr_gpr_iu_gpr_15__25_), .Y(_6118_) );
	OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf4), .B(_6092__bF_buf4), .C(_6118_), .Y(_1845_) );
	OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6026__bF_buf6), .C(csr_gpr_iu_gpr_15__26_), .Y(_6119_) );
	OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf4), .B(_6092__bF_buf3), .C(_6119_), .Y(_1846_) );
	OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6026__bF_buf5), .C(csr_gpr_iu_gpr_15__27_), .Y(_6120_) );
	OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf4), .B(_6092__bF_buf2), .C(_6120_), .Y(_1847_) );
	OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6026__bF_buf4), .C(csr_gpr_iu_gpr_15__28_), .Y(_6121_) );
	OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf4), .B(_6092__bF_buf1), .C(_6121_), .Y(_1848_) );
	OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6026__bF_buf3), .C(csr_gpr_iu_gpr_15__29_), .Y(_6122_) );
	OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf4), .B(_6092__bF_buf0), .C(_6122_), .Y(_1849_) );
	OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6026__bF_buf2), .C(csr_gpr_iu_gpr_15__30_), .Y(_6123_) );
	OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_6092__bF_buf4), .C(_6123_), .Y(_1850_) );
	OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6026__bF_buf1), .C(csr_gpr_iu_gpr_15__31_), .Y(_6124_) );
	OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf4), .B(_6092__bF_buf3), .C(_6124_), .Y(_1851_) );
	NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_2993__bF_buf0), .B(_2484__bF_buf12), .Y(_6125_) );
	NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_0_), .B(_2995__bF_buf6), .C(_2473__bF_buf5), .Y(_6126_) );
	OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_6125__bF_buf4), .C(_6126_), .Y(_1852_) );
	NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_1_), .B(_2995__bF_buf5), .C(_2473__bF_buf4), .Y(_6127_) );
	OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_6125__bF_buf3), .C(_6127_), .Y(_1853_) );
	NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_2_), .B(_2995__bF_buf4), .C(_2473__bF_buf3), .Y(_6128_) );
	OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_6125__bF_buf2), .C(_6128_), .Y(_1854_) );
	NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_3_), .B(_2995__bF_buf3), .C(_2473__bF_buf2), .Y(_6129_) );
	OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_6125__bF_buf1), .C(_6129_), .Y(_1855_) );
	NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_4_), .B(_2995__bF_buf2), .C(_2473__bF_buf1), .Y(_6130_) );
	OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(_6125__bF_buf0), .C(_6130_), .Y(_1856_) );
	NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_5_), .B(_2995__bF_buf1), .C(_2473__bF_buf0), .Y(_6131_) );
	OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_6125__bF_buf4), .C(_6131_), .Y(_1857_) );
	NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_6_), .B(_2995__bF_buf0), .C(_2473__bF_buf7), .Y(_6132_) );
	OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_6125__bF_buf3), .C(_6132_), .Y(_1858_) );
	NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_7_), .B(_2995__bF_buf8), .C(_2473__bF_buf6), .Y(_6133_) );
	OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_6125__bF_buf2), .C(_6133_), .Y(_1859_) );
	NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_8_), .B(_2995__bF_buf7), .C(_2473__bF_buf5), .Y(_6134_) );
	OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_6125__bF_buf1), .C(_6134_), .Y(_1860_) );
	NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_9_), .B(_2995__bF_buf6), .C(_2473__bF_buf4), .Y(_6135_) );
	OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(_6125__bF_buf0), .C(_6135_), .Y(_1861_) );
	NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_10_), .B(_2995__bF_buf5), .C(_2473__bF_buf3), .Y(_6136_) );
	OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_6125__bF_buf4), .C(_6136_), .Y(_1862_) );
	NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_11_), .B(_2995__bF_buf4), .C(_2473__bF_buf2), .Y(_6137_) );
	OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_3770_), .B(_6125__bF_buf3), .C(_6137_), .Y(_1863_) );
	NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_12_), .B(_2995__bF_buf3), .C(_2473__bF_buf1), .Y(_6138_) );
	OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_3794_), .B(_6125__bF_buf2), .C(_6138_), .Y(_1864_) );
	NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_13_), .B(_2995__bF_buf2), .C(_2473__bF_buf0), .Y(_6139_) );
	OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_3880_), .B(_6125__bF_buf1), .C(_6139_), .Y(_1865_) );
	NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_14_), .B(_2995__bF_buf1), .C(_2473__bF_buf7), .Y(_6140_) );
	OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_6125__bF_buf0), .C(_6140_), .Y(_1866_) );
	NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_15_), .B(_2995__bF_buf0), .C(_2473__bF_buf6), .Y(_6141_) );
	OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_6125__bF_buf4), .C(_6141_), .Y(_1867_) );
	NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_16_), .B(_2995__bF_buf8), .C(_2473__bF_buf5), .Y(_6142_) );
	OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_6125__bF_buf3), .C(_6142_), .Y(_1868_) );
	NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_17_), .B(_2995__bF_buf7), .C(_2473__bF_buf4), .Y(_6143_) );
	OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_6125__bF_buf2), .C(_6143_), .Y(_1869_) );
	NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_18_), .B(_2995__bF_buf6), .C(_2473__bF_buf3), .Y(_6144_) );
	OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(_6125__bF_buf1), .C(_6144_), .Y(_1870_) );
	NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_19_), .B(_2995__bF_buf5), .C(_2473__bF_buf2), .Y(_6145_) );
	OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_4210_), .B(_6125__bF_buf0), .C(_6145_), .Y(_1871_) );
	NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_20_), .B(_2995__bF_buf4), .C(_2473__bF_buf1), .Y(_6146_) );
	OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .B(_6125__bF_buf4), .C(_6146_), .Y(_1872_) );
	NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_21_), .B(_2995__bF_buf3), .C(_2473__bF_buf0), .Y(_6147_) );
	OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_4320_), .B(_6125__bF_buf3), .C(_6147_), .Y(_1873_) );
	NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_22_), .B(_2995__bF_buf2), .C(_2473__bF_buf7), .Y(_6148_) );
	OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_4375_), .B(_6125__bF_buf2), .C(_6148_), .Y(_1874_) );
	NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_23_), .B(_2995__bF_buf1), .C(_2473__bF_buf6), .Y(_6149_) );
	OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_6125__bF_buf1), .C(_6149_), .Y(_1875_) );
	NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_24_), .B(_2995__bF_buf0), .C(_2473__bF_buf5), .Y(_6150_) );
	OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_4454_), .B(_6125__bF_buf0), .C(_6150_), .Y(_1876_) );
	NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_25_), .B(_2995__bF_buf8), .C(_2473__bF_buf4), .Y(_6151_) );
	OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_4509_), .B(_6125__bF_buf4), .C(_6151_), .Y(_1877_) );
	NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_26_), .B(_2995__bF_buf7), .C(_2473__bF_buf3), .Y(_6152_) );
	OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_6125__bF_buf3), .C(_6152_), .Y(_1878_) );
	NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_27_), .B(_2995__bF_buf6), .C(_2473__bF_buf2), .Y(_6153_) );
	OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_4650_), .B(_6125__bF_buf2), .C(_6153_), .Y(_1879_) );
	NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_28_), .B(_2995__bF_buf5), .C(_2473__bF_buf1), .Y(_6154_) );
	OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .B(_6125__bF_buf1), .C(_6154_), .Y(_1880_) );
	NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_29_), .B(_2995__bF_buf4), .C(_2473__bF_buf0), .Y(_6155_) );
	OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_6125__bF_buf0), .C(_6155_), .Y(_1881_) );
	NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_30_), .B(_2995__bF_buf3), .C(_2473__bF_buf7), .Y(_6156_) );
	OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_6125__bF_buf4), .C(_6156_), .Y(_1882_) );
	NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_data_gpr_31_), .B(_2995__bF_buf2), .C(_2473__bF_buf6), .Y(_6157_) );
	OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_4870_), .B(_6125__bF_buf3), .C(_6157_), .Y(_1883_) );
	NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .B(_2486_), .Y(_6158_) );
	NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_6158_), .C(_2694__bF_buf5), .Y(_6159_) );
	NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_6158_), .Y(_6160_) );
	OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_0__0_), .Y(_6161_) );
	OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf3), .B(_6159__bF_buf4), .C(_6161_), .Y(_1884_) );
	OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_0__1_), .Y(_6162_) );
	OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf3), .B(_6159__bF_buf3), .C(_6162_), .Y(_1885_) );
	OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_0__2_), .Y(_6163_) );
	OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf3), .B(_6159__bF_buf2), .C(_6163_), .Y(_1886_) );
	OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_0__3_), .Y(_6164_) );
	OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf3), .B(_6159__bF_buf1), .C(_6164_), .Y(_1887_) );
	OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_0__4_), .Y(_6165_) );
	OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf3), .B(_6159__bF_buf0), .C(_6165_), .Y(_1888_) );
	OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_0__5_), .Y(_6166_) );
	OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf3), .B(_6159__bF_buf4), .C(_6166_), .Y(_1889_) );
	OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_0__6_), .Y(_6167_) );
	OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf3), .B(_6159__bF_buf3), .C(_6167_), .Y(_1890_) );
	OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_0__7_), .Y(_6168_) );
	OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf3), .B(_6159__bF_buf2), .C(_6168_), .Y(_1891_) );
	OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_0__8_), .Y(_6169_) );
	OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf3), .B(_6159__bF_buf1), .C(_6169_), .Y(_1892_) );
	OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_0__9_), .Y(_6170_) );
	OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf3), .B(_6159__bF_buf0), .C(_6170_), .Y(_1893_) );
	OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_0__10_), .Y(_6171_) );
	OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf3), .B(_6159__bF_buf4), .C(_6171_), .Y(_1894_) );
	OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_0__11_), .Y(_6172_) );
	OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf3), .B(_6159__bF_buf3), .C(_6172_), .Y(_1895_) );
	OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_0__12_), .Y(_6173_) );
	OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf3), .B(_6159__bF_buf2), .C(_6173_), .Y(_1896_) );
	OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_0__13_), .Y(_6174_) );
	OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf3), .B(_6159__bF_buf1), .C(_6174_), .Y(_1897_) );
	OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_0__14_), .Y(_6175_) );
	OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf3), .B(_6159__bF_buf0), .C(_6175_), .Y(_1898_) );
	OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_0__15_), .Y(_6176_) );
	OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf3), .B(_6159__bF_buf4), .C(_6176_), .Y(_1899_) );
	OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_0__16_), .Y(_6177_) );
	OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf3), .B(_6159__bF_buf3), .C(_6177_), .Y(_1900_) );
	OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_0__17_), .Y(_6178_) );
	OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf3), .B(_6159__bF_buf2), .C(_6178_), .Y(_1901_) );
	OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_0__18_), .Y(_6179_) );
	OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf3), .B(_6159__bF_buf1), .C(_6179_), .Y(_1902_) );
	OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_0__19_), .Y(_6180_) );
	OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf3), .B(_6159__bF_buf0), .C(_6180_), .Y(_1903_) );
	OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_0__20_), .Y(_6181_) );
	OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf3), .B(_6159__bF_buf4), .C(_6181_), .Y(_1904_) );
	OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_0__21_), .Y(_6182_) );
	OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf3), .B(_6159__bF_buf3), .C(_6182_), .Y(_1905_) );
	OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_0__22_), .Y(_6183_) );
	OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf3), .B(_6159__bF_buf2), .C(_6183_), .Y(_1906_) );
	OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_0__23_), .Y(_6184_) );
	OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf3), .B(_6159__bF_buf1), .C(_6184_), .Y(_1907_) );
	OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_0__24_), .Y(_6185_) );
	OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf3), .B(_6159__bF_buf0), .C(_6185_), .Y(_1908_) );
	OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_0__25_), .Y(_6186_) );
	OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf3), .B(_6159__bF_buf4), .C(_6186_), .Y(_1909_) );
	OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_0__26_), .Y(_6187_) );
	OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf3), .B(_6159__bF_buf3), .C(_6187_), .Y(_1910_) );
	OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_0__27_), .Y(_6188_) );
	OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf3), .B(_6159__bF_buf2), .C(_6188_), .Y(_1911_) );
	OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_0__28_), .Y(_6189_) );
	OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf3), .B(_6159__bF_buf1), .C(_6189_), .Y(_1912_) );
	OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_0__29_), .Y(_6190_) );
	OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf3), .B(_6159__bF_buf0), .C(_6190_), .Y(_1913_) );
	OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_0__30_), .Y(_6191_) );
	OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_6159__bF_buf4), .C(_6191_), .Y(_1914_) );
	OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_0__31_), .Y(_6192_) );
	OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf3), .B(_6159__bF_buf3), .C(_6192_), .Y(_1915_) );
	NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_6158_), .C(_2473__bF_buf5), .Y(_6193_) );
	OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_1__0_), .Y(_6194_) );
	OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf2), .B(_6193__bF_buf4), .C(_6194_), .Y(_1916_) );
	OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_1__1_), .Y(_6195_) );
	OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf2), .B(_6193__bF_buf3), .C(_6195_), .Y(_1917_) );
	OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_1__2_), .Y(_6196_) );
	OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf2), .B(_6193__bF_buf2), .C(_6196_), .Y(_1918_) );
	OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_1__3_), .Y(_6197_) );
	OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf2), .B(_6193__bF_buf1), .C(_6197_), .Y(_1919_) );
	OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_1__4_), .Y(_6198_) );
	OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf2), .B(_6193__bF_buf0), .C(_6198_), .Y(_1920_) );
	OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_1__5_), .Y(_6199_) );
	OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf2), .B(_6193__bF_buf4), .C(_6199_), .Y(_1921_) );
	OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_1__6_), .Y(_6200_) );
	OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf2), .B(_6193__bF_buf3), .C(_6200_), .Y(_1922_) );
	OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_1__7_), .Y(_6201_) );
	OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf2), .B(_6193__bF_buf2), .C(_6201_), .Y(_1923_) );
	OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_1__8_), .Y(_6202_) );
	OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf2), .B(_6193__bF_buf1), .C(_6202_), .Y(_1924_) );
	OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_1__9_), .Y(_6203_) );
	OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf2), .B(_6193__bF_buf0), .C(_6203_), .Y(_1925_) );
	OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_1__10_), .Y(_6204_) );
	OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf2), .B(_6193__bF_buf4), .C(_6204_), .Y(_1926_) );
	OAI21X1 OAI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_1__11_), .Y(_6205_) );
	OAI21X1 OAI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf2), .B(_6193__bF_buf3), .C(_6205_), .Y(_1927_) );
	OAI21X1 OAI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_1__12_), .Y(_6206_) );
	OAI21X1 OAI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf2), .B(_6193__bF_buf2), .C(_6206_), .Y(_1928_) );
	OAI21X1 OAI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_1__13_), .Y(_6207_) );
	OAI21X1 OAI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf2), .B(_6193__bF_buf1), .C(_6207_), .Y(_1929_) );
	OAI21X1 OAI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_1__14_), .Y(_6208_) );
	OAI21X1 OAI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf2), .B(_6193__bF_buf0), .C(_6208_), .Y(_1930_) );
	OAI21X1 OAI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_1__15_), .Y(_6209_) );
	OAI21X1 OAI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf2), .B(_6193__bF_buf4), .C(_6209_), .Y(_1931_) );
	OAI21X1 OAI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_1__16_), .Y(_6210_) );
	OAI21X1 OAI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf2), .B(_6193__bF_buf3), .C(_6210_), .Y(_1932_) );
	OAI21X1 OAI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_1__17_), .Y(_6211_) );
	OAI21X1 OAI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf2), .B(_6193__bF_buf2), .C(_6211_), .Y(_1933_) );
	OAI21X1 OAI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_1__18_), .Y(_6212_) );
	OAI21X1 OAI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf2), .B(_6193__bF_buf1), .C(_6212_), .Y(_1934_) );
	OAI21X1 OAI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_1__19_), .Y(_6213_) );
	OAI21X1 OAI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf2), .B(_6193__bF_buf0), .C(_6213_), .Y(_1935_) );
	OAI21X1 OAI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_1__20_), .Y(_6214_) );
	OAI21X1 OAI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf2), .B(_6193__bF_buf4), .C(_6214_), .Y(_1936_) );
	OAI21X1 OAI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_1__21_), .Y(_6215_) );
	OAI21X1 OAI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf2), .B(_6193__bF_buf3), .C(_6215_), .Y(_1937_) );
	OAI21X1 OAI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_1__22_), .Y(_6216_) );
	OAI21X1 OAI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf2), .B(_6193__bF_buf2), .C(_6216_), .Y(_1938_) );
	OAI21X1 OAI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_1__23_), .Y(_6217_) );
	OAI21X1 OAI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf2), .B(_6193__bF_buf1), .C(_6217_), .Y(_1939_) );
	OAI21X1 OAI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_1__24_), .Y(_6218_) );
	OAI21X1 OAI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf2), .B(_6193__bF_buf0), .C(_6218_), .Y(_1940_) );
	OAI21X1 OAI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_1__25_), .Y(_6219_) );
	OAI21X1 OAI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf2), .B(_6193__bF_buf4), .C(_6219_), .Y(_1941_) );
	OAI21X1 OAI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_1__26_), .Y(_6220_) );
	OAI21X1 OAI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf2), .B(_6193__bF_buf3), .C(_6220_), .Y(_1942_) );
	OAI21X1 OAI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_1__27_), .Y(_6221_) );
	OAI21X1 OAI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf2), .B(_6193__bF_buf2), .C(_6221_), .Y(_1943_) );
	OAI21X1 OAI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_1__28_), .Y(_6222_) );
	OAI21X1 OAI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf2), .B(_6193__bF_buf1), .C(_6222_), .Y(_1944_) );
	OAI21X1 OAI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_1__29_), .Y(_6223_) );
	OAI21X1 OAI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf2), .B(_6193__bF_buf0), .C(_6223_), .Y(_1945_) );
	OAI21X1 OAI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_1__30_), .Y(_6224_) );
	OAI21X1 OAI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_6193__bF_buf4), .C(_6224_), .Y(_1946_) );
	OAI21X1 OAI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_1__31_), .Y(_6225_) );
	OAI21X1 OAI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf2), .B(_6193__bF_buf3), .C(_6225_), .Y(_1947_) );
	NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_6158_), .C(_2588__bF_buf4), .Y(_6226_) );
	OAI21X1 OAI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_2__0_), .Y(_6227_) );
	OAI21X1 OAI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf1), .B(_6226__bF_buf4), .C(_6227_), .Y(_1948_) );
	OAI21X1 OAI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_2__1_), .Y(_6228_) );
	OAI21X1 OAI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf1), .B(_6226__bF_buf3), .C(_6228_), .Y(_1949_) );
	OAI21X1 OAI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_2__2_), .Y(_6229_) );
	OAI21X1 OAI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf1), .B(_6226__bF_buf2), .C(_6229_), .Y(_1950_) );
	OAI21X1 OAI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_2__3_), .Y(_6230_) );
	OAI21X1 OAI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf1), .B(_6226__bF_buf1), .C(_6230_), .Y(_1951_) );
	OAI21X1 OAI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_2__4_), .Y(_6231_) );
	OAI21X1 OAI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf1), .B(_6226__bF_buf0), .C(_6231_), .Y(_1952_) );
	OAI21X1 OAI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_2__5_), .Y(_6232_) );
	OAI21X1 OAI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf1), .B(_6226__bF_buf4), .C(_6232_), .Y(_1953_) );
	OAI21X1 OAI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_2__6_), .Y(_6233_) );
	OAI21X1 OAI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf1), .B(_6226__bF_buf3), .C(_6233_), .Y(_1954_) );
	OAI21X1 OAI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_2__7_), .Y(_6234_) );
	OAI21X1 OAI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf1), .B(_6226__bF_buf2), .C(_6234_), .Y(_1955_) );
	OAI21X1 OAI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_2__8_), .Y(_6235_) );
	OAI21X1 OAI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf1), .B(_6226__bF_buf1), .C(_6235_), .Y(_1956_) );
	OAI21X1 OAI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_2__9_), .Y(_6236_) );
	OAI21X1 OAI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf1), .B(_6226__bF_buf0), .C(_6236_), .Y(_1957_) );
	OAI21X1 OAI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_2__10_), .Y(_6237_) );
	OAI21X1 OAI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf1), .B(_6226__bF_buf4), .C(_6237_), .Y(_1958_) );
	OAI21X1 OAI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_2__11_), .Y(_6238_) );
	OAI21X1 OAI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf1), .B(_6226__bF_buf3), .C(_6238_), .Y(_1959_) );
	OAI21X1 OAI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_2__12_), .Y(_6239_) );
	OAI21X1 OAI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf1), .B(_6226__bF_buf2), .C(_6239_), .Y(_1960_) );
	OAI21X1 OAI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_2__13_), .Y(_6240_) );
	OAI21X1 OAI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf1), .B(_6226__bF_buf1), .C(_6240_), .Y(_1961_) );
	OAI21X1 OAI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_2__14_), .Y(_6241_) );
	OAI21X1 OAI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf1), .B(_6226__bF_buf0), .C(_6241_), .Y(_1962_) );
	OAI21X1 OAI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_2__15_), .Y(_6242_) );
	OAI21X1 OAI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf1), .B(_6226__bF_buf4), .C(_6242_), .Y(_1963_) );
	OAI21X1 OAI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_2__16_), .Y(_6243_) );
	OAI21X1 OAI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf1), .B(_6226__bF_buf3), .C(_6243_), .Y(_1964_) );
	OAI21X1 OAI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_2__17_), .Y(_6244_) );
	OAI21X1 OAI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf1), .B(_6226__bF_buf2), .C(_6244_), .Y(_1965_) );
	OAI21X1 OAI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_2__18_), .Y(_6245_) );
	OAI21X1 OAI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf1), .B(_6226__bF_buf1), .C(_6245_), .Y(_1966_) );
	OAI21X1 OAI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_2__19_), .Y(_6246_) );
	OAI21X1 OAI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf1), .B(_6226__bF_buf0), .C(_6246_), .Y(_1967_) );
	OAI21X1 OAI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_2__20_), .Y(_6247_) );
	OAI21X1 OAI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf1), .B(_6226__bF_buf4), .C(_6247_), .Y(_1968_) );
	OAI21X1 OAI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_2__21_), .Y(_6248_) );
	OAI21X1 OAI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf1), .B(_6226__bF_buf3), .C(_6248_), .Y(_1969_) );
	OAI21X1 OAI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_2__22_), .Y(_6249_) );
	OAI21X1 OAI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf1), .B(_6226__bF_buf2), .C(_6249_), .Y(_1970_) );
	OAI21X1 OAI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_2__23_), .Y(_6250_) );
	OAI21X1 OAI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf1), .B(_6226__bF_buf1), .C(_6250_), .Y(_1971_) );
	OAI21X1 OAI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_2__24_), .Y(_6251_) );
	OAI21X1 OAI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf1), .B(_6226__bF_buf0), .C(_6251_), .Y(_1972_) );
	OAI21X1 OAI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_2__25_), .Y(_6252_) );
	OAI21X1 OAI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf1), .B(_6226__bF_buf4), .C(_6252_), .Y(_1973_) );
	OAI21X1 OAI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_2__26_), .Y(_6253_) );
	OAI21X1 OAI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf1), .B(_6226__bF_buf3), .C(_6253_), .Y(_1974_) );
	OAI21X1 OAI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_2__27_), .Y(_6254_) );
	OAI21X1 OAI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf1), .B(_6226__bF_buf2), .C(_6254_), .Y(_1975_) );
	OAI21X1 OAI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_2__28_), .Y(_6255_) );
	OAI21X1 OAI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf1), .B(_6226__bF_buf1), .C(_6255_), .Y(_1976_) );
	OAI21X1 OAI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_2__29_), .Y(_6256_) );
	OAI21X1 OAI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf1), .B(_6226__bF_buf0), .C(_6256_), .Y(_1977_) );
	OAI21X1 OAI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_2__30_), .Y(_6257_) );
	OAI21X1 OAI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_6226__bF_buf4), .C(_6257_), .Y(_1978_) );
	OAI21X1 OAI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_2__31_), .Y(_6258_) );
	OAI21X1 OAI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf1), .B(_6226__bF_buf3), .C(_6258_), .Y(_1979_) );
	NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_6158_), .C(_2623_), .Y(_6259_) );
	OAI21X1 OAI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_3__0_), .Y(_6260_) );
	OAI21X1 OAI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf0), .B(_6259__bF_buf4), .C(_6260_), .Y(_1980_) );
	OAI21X1 OAI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_3__1_), .Y(_6261_) );
	OAI21X1 OAI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf0), .B(_6259__bF_buf3), .C(_6261_), .Y(_1981_) );
	OAI21X1 OAI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_3__2_), .Y(_6262_) );
	OAI21X1 OAI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf0), .B(_6259__bF_buf2), .C(_6262_), .Y(_1982_) );
	OAI21X1 OAI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_3__3_), .Y(_6263_) );
	OAI21X1 OAI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf0), .B(_6259__bF_buf1), .C(_6263_), .Y(_1983_) );
	OAI21X1 OAI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_3__4_), .Y(_6264_) );
	OAI21X1 OAI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf0), .B(_6259__bF_buf0), .C(_6264_), .Y(_1984_) );
	OAI21X1 OAI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_3__5_), .Y(_6265_) );
	OAI21X1 OAI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf0), .B(_6259__bF_buf4), .C(_6265_), .Y(_1985_) );
	OAI21X1 OAI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_3__6_), .Y(_6266_) );
	OAI21X1 OAI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf0), .B(_6259__bF_buf3), .C(_6266_), .Y(_1986_) );
	OAI21X1 OAI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_3__7_), .Y(_6267_) );
	OAI21X1 OAI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf0), .B(_6259__bF_buf2), .C(_6267_), .Y(_1987_) );
	OAI21X1 OAI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_3__8_), .Y(_6268_) );
	OAI21X1 OAI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf0), .B(_6259__bF_buf1), .C(_6268_), .Y(_1988_) );
	OAI21X1 OAI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_3__9_), .Y(_6269_) );
	OAI21X1 OAI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf0), .B(_6259__bF_buf0), .C(_6269_), .Y(_1989_) );
	OAI21X1 OAI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_3__10_), .Y(_6270_) );
	OAI21X1 OAI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf0), .B(_6259__bF_buf4), .C(_6270_), .Y(_1990_) );
	OAI21X1 OAI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_3__11_), .Y(_6271_) );
	OAI21X1 OAI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf0), .B(_6259__bF_buf3), .C(_6271_), .Y(_1991_) );
	OAI21X1 OAI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_3__12_), .Y(_6272_) );
	OAI21X1 OAI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf0), .B(_6259__bF_buf2), .C(_6272_), .Y(_1992_) );
	OAI21X1 OAI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_3__13_), .Y(_6273_) );
	OAI21X1 OAI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf0), .B(_6259__bF_buf1), .C(_6273_), .Y(_1993_) );
	OAI21X1 OAI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_3__14_), .Y(_6274_) );
	OAI21X1 OAI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf0), .B(_6259__bF_buf0), .C(_6274_), .Y(_1994_) );
	OAI21X1 OAI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_3__15_), .Y(_6275_) );
	OAI21X1 OAI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf0), .B(_6259__bF_buf4), .C(_6275_), .Y(_1995_) );
	OAI21X1 OAI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_3__16_), .Y(_6276_) );
	OAI21X1 OAI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf0), .B(_6259__bF_buf3), .C(_6276_), .Y(_1996_) );
	OAI21X1 OAI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_3__17_), .Y(_6277_) );
	OAI21X1 OAI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf0), .B(_6259__bF_buf2), .C(_6277_), .Y(_1997_) );
	OAI21X1 OAI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_3__18_), .Y(_6278_) );
	OAI21X1 OAI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf0), .B(_6259__bF_buf1), .C(_6278_), .Y(_1998_) );
	OAI21X1 OAI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_3__19_), .Y(_6279_) );
	OAI21X1 OAI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf0), .B(_6259__bF_buf0), .C(_6279_), .Y(_1999_) );
	OAI21X1 OAI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_3__20_), .Y(_6280_) );
	OAI21X1 OAI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf0), .B(_6259__bF_buf4), .C(_6280_), .Y(_2000_) );
	OAI21X1 OAI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6160__bF_buf3), .C(csr_gpr_iu_gpr_3__21_), .Y(_6281_) );
	OAI21X1 OAI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf0), .B(_6259__bF_buf3), .C(_6281_), .Y(_2001_) );
	OAI21X1 OAI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6160__bF_buf2), .C(csr_gpr_iu_gpr_3__22_), .Y(_6282_) );
	OAI21X1 OAI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf0), .B(_6259__bF_buf2), .C(_6282_), .Y(_2002_) );
	OAI21X1 OAI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6160__bF_buf1), .C(csr_gpr_iu_gpr_3__23_), .Y(_6283_) );
	OAI21X1 OAI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf0), .B(_6259__bF_buf1), .C(_6283_), .Y(_2003_) );
	OAI21X1 OAI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6160__bF_buf0), .C(csr_gpr_iu_gpr_3__24_), .Y(_6284_) );
	OAI21X1 OAI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf0), .B(_6259__bF_buf0), .C(_6284_), .Y(_2004_) );
	OAI21X1 OAI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6160__bF_buf10), .C(csr_gpr_iu_gpr_3__25_), .Y(_6285_) );
	OAI21X1 OAI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf0), .B(_6259__bF_buf4), .C(_6285_), .Y(_2005_) );
	OAI21X1 OAI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6160__bF_buf9), .C(csr_gpr_iu_gpr_3__26_), .Y(_6286_) );
	OAI21X1 OAI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf0), .B(_6259__bF_buf3), .C(_6286_), .Y(_2006_) );
	OAI21X1 OAI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6160__bF_buf8), .C(csr_gpr_iu_gpr_3__27_), .Y(_6287_) );
	OAI21X1 OAI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf0), .B(_6259__bF_buf2), .C(_6287_), .Y(_2007_) );
	OAI21X1 OAI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6160__bF_buf7), .C(csr_gpr_iu_gpr_3__28_), .Y(_6288_) );
	OAI21X1 OAI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf0), .B(_6259__bF_buf1), .C(_6288_), .Y(_2008_) );
	OAI21X1 OAI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6160__bF_buf6), .C(csr_gpr_iu_gpr_3__29_), .Y(_6289_) );
	OAI21X1 OAI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf0), .B(_6259__bF_buf0), .C(_6289_), .Y(_2009_) );
	OAI21X1 OAI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6160__bF_buf5), .C(csr_gpr_iu_gpr_3__30_), .Y(_6290_) );
	OAI21X1 OAI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_6259__bF_buf4), .C(_6290_), .Y(_2010_) );
	OAI21X1 OAI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6160__bF_buf4), .C(csr_gpr_iu_gpr_3__31_), .Y(_6291_) );
	OAI21X1 OAI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf0), .B(_6259__bF_buf3), .C(_6291_), .Y(_2011_) );
	NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_6158_), .C(_2694__bF_buf4), .Y(_6292_) );
	NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_6158_), .Y(_6293_) );
	OAI21X1 OAI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_4__0_), .Y(_6294_) );
	OAI21X1 OAI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf4), .B(_6292__bF_buf4), .C(_6294_), .Y(_2012_) );
	OAI21X1 OAI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_4__1_), .Y(_6295_) );
	OAI21X1 OAI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf4), .B(_6292__bF_buf3), .C(_6295_), .Y(_2013_) );
	OAI21X1 OAI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_4__2_), .Y(_6296_) );
	OAI21X1 OAI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf4), .B(_6292__bF_buf2), .C(_6296_), .Y(_2014_) );
	OAI21X1 OAI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_4__3_), .Y(_6297_) );
	OAI21X1 OAI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf4), .B(_6292__bF_buf1), .C(_6297_), .Y(_2015_) );
	OAI21X1 OAI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_4__4_), .Y(_6298_) );
	OAI21X1 OAI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf4), .B(_6292__bF_buf0), .C(_6298_), .Y(_2016_) );
	OAI21X1 OAI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_4__5_), .Y(_6299_) );
	OAI21X1 OAI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf4), .B(_6292__bF_buf4), .C(_6299_), .Y(_2017_) );
	OAI21X1 OAI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_4__6_), .Y(_6300_) );
	OAI21X1 OAI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf4), .B(_6292__bF_buf3), .C(_6300_), .Y(_2018_) );
	OAI21X1 OAI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_4__7_), .Y(_6301_) );
	OAI21X1 OAI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf4), .B(_6292__bF_buf2), .C(_6301_), .Y(_2019_) );
	OAI21X1 OAI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_4__8_), .Y(_6302_) );
	OAI21X1 OAI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf4), .B(_6292__bF_buf1), .C(_6302_), .Y(_2020_) );
	OAI21X1 OAI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_4__9_), .Y(_6303_) );
	OAI21X1 OAI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf4), .B(_6292__bF_buf0), .C(_6303_), .Y(_2021_) );
	OAI21X1 OAI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_4__10_), .Y(_6304_) );
	OAI21X1 OAI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf4), .B(_6292__bF_buf4), .C(_6304_), .Y(_2022_) );
	OAI21X1 OAI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_4__11_), .Y(_6305_) );
	OAI21X1 OAI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf4), .B(_6292__bF_buf3), .C(_6305_), .Y(_2023_) );
	OAI21X1 OAI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_4__12_), .Y(_6306_) );
	OAI21X1 OAI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf4), .B(_6292__bF_buf2), .C(_6306_), .Y(_2024_) );
	OAI21X1 OAI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_4__13_), .Y(_6307_) );
	OAI21X1 OAI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf4), .B(_6292__bF_buf1), .C(_6307_), .Y(_2025_) );
	OAI21X1 OAI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_4__14_), .Y(_6308_) );
	OAI21X1 OAI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf4), .B(_6292__bF_buf0), .C(_6308_), .Y(_2026_) );
	OAI21X1 OAI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_4__15_), .Y(_6309_) );
	OAI21X1 OAI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf4), .B(_6292__bF_buf4), .C(_6309_), .Y(_2027_) );
	OAI21X1 OAI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_4__16_), .Y(_6310_) );
	OAI21X1 OAI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf4), .B(_6292__bF_buf3), .C(_6310_), .Y(_2028_) );
	OAI21X1 OAI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_4__17_), .Y(_6311_) );
	OAI21X1 OAI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf4), .B(_6292__bF_buf2), .C(_6311_), .Y(_2029_) );
	OAI21X1 OAI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_4__18_), .Y(_6312_) );
	OAI21X1 OAI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf4), .B(_6292__bF_buf1), .C(_6312_), .Y(_2030_) );
	OAI21X1 OAI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf12), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_4__19_), .Y(_6313_) );
	OAI21X1 OAI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf4), .B(_6292__bF_buf0), .C(_6313_), .Y(_2031_) );
	OAI21X1 OAI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf11), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_4__20_), .Y(_6314_) );
	OAI21X1 OAI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf4), .B(_6292__bF_buf4), .C(_6314_), .Y(_2032_) );
	OAI21X1 OAI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf10), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_4__21_), .Y(_6315_) );
	OAI21X1 OAI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf4), .B(_6292__bF_buf3), .C(_6315_), .Y(_2033_) );
	OAI21X1 OAI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf9), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_4__22_), .Y(_6316_) );
	OAI21X1 OAI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf4), .B(_6292__bF_buf2), .C(_6316_), .Y(_2034_) );
	OAI21X1 OAI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf8), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_4__23_), .Y(_6317_) );
	OAI21X1 OAI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf4), .B(_6292__bF_buf1), .C(_6317_), .Y(_2035_) );
	OAI21X1 OAI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf7), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_4__24_), .Y(_6318_) );
	OAI21X1 OAI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf4), .B(_6292__bF_buf0), .C(_6318_), .Y(_2036_) );
	OAI21X1 OAI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf6), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_4__25_), .Y(_6319_) );
	OAI21X1 OAI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf4), .B(_6292__bF_buf4), .C(_6319_), .Y(_2037_) );
	OAI21X1 OAI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf5), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_4__26_), .Y(_6320_) );
	OAI21X1 OAI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf4), .B(_6292__bF_buf3), .C(_6320_), .Y(_2038_) );
	OAI21X1 OAI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf4), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_4__27_), .Y(_6321_) );
	OAI21X1 OAI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf4), .B(_6292__bF_buf2), .C(_6321_), .Y(_2039_) );
	OAI21X1 OAI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf3), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_4__28_), .Y(_6322_) );
	OAI21X1 OAI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf4), .B(_6292__bF_buf1), .C(_6322_), .Y(_2040_) );
	OAI21X1 OAI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf2), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_4__29_), .Y(_6323_) );
	OAI21X1 OAI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf4), .B(_6292__bF_buf0), .C(_6323_), .Y(_2041_) );
	OAI21X1 OAI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf1), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_4__30_), .Y(_6324_) );
	OAI21X1 OAI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_6292__bF_buf4), .C(_6324_), .Y(_2042_) );
	OAI21X1 OAI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_2696__bF_buf0), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_4__31_), .Y(_6325_) );
	OAI21X1 OAI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf4), .B(_6292__bF_buf3), .C(_6325_), .Y(_2043_) );
	NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_6158_), .C(_2473__bF_buf4), .Y(_6326_) );
	OAI21X1 OAI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_5__0_), .Y(_6327_) );
	OAI21X1 OAI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf3), .B(_6326__bF_buf4), .C(_6327_), .Y(_2044_) );
	OAI21X1 OAI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_5__1_), .Y(_6328_) );
	OAI21X1 OAI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf3), .B(_6326__bF_buf3), .C(_6328_), .Y(_2045_) );
	OAI21X1 OAI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_5__2_), .Y(_6329_) );
	OAI21X1 OAI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf3), .B(_6326__bF_buf2), .C(_6329_), .Y(_2046_) );
	OAI21X1 OAI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_5__3_), .Y(_6330_) );
	OAI21X1 OAI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf3), .B(_6326__bF_buf1), .C(_6330_), .Y(_2047_) );
	OAI21X1 OAI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_5__4_), .Y(_6331_) );
	OAI21X1 OAI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf3), .B(_6326__bF_buf0), .C(_6331_), .Y(_2048_) );
	OAI21X1 OAI21X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_5__5_), .Y(_6332_) );
	OAI21X1 OAI21X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf3), .B(_6326__bF_buf4), .C(_6332_), .Y(_2049_) );
	OAI21X1 OAI21X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_5__6_), .Y(_6333_) );
	OAI21X1 OAI21X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf3), .B(_6326__bF_buf3), .C(_6333_), .Y(_2050_) );
	OAI21X1 OAI21X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_5__7_), .Y(_6334_) );
	OAI21X1 OAI21X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf3), .B(_6326__bF_buf2), .C(_6334_), .Y(_2051_) );
	OAI21X1 OAI21X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_5__8_), .Y(_6335_) );
	OAI21X1 OAI21X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf3), .B(_6326__bF_buf1), .C(_6335_), .Y(_2052_) );
	OAI21X1 OAI21X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_5__9_), .Y(_6336_) );
	OAI21X1 OAI21X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf3), .B(_6326__bF_buf0), .C(_6336_), .Y(_2053_) );
	OAI21X1 OAI21X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_5__10_), .Y(_6337_) );
	OAI21X1 OAI21X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf3), .B(_6326__bF_buf4), .C(_6337_), .Y(_2054_) );
	OAI21X1 OAI21X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_5__11_), .Y(_6338_) );
	OAI21X1 OAI21X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf3), .B(_6326__bF_buf3), .C(_6338_), .Y(_2055_) );
	OAI21X1 OAI21X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_5__12_), .Y(_6339_) );
	OAI21X1 OAI21X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf3), .B(_6326__bF_buf2), .C(_6339_), .Y(_2056_) );
	OAI21X1 OAI21X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_5__13_), .Y(_6340_) );
	OAI21X1 OAI21X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf3), .B(_6326__bF_buf1), .C(_6340_), .Y(_2057_) );
	OAI21X1 OAI21X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_5__14_), .Y(_6341_) );
	OAI21X1 OAI21X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf3), .B(_6326__bF_buf0), .C(_6341_), .Y(_2058_) );
	OAI21X1 OAI21X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_5__15_), .Y(_6342_) );
	OAI21X1 OAI21X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf3), .B(_6326__bF_buf4), .C(_6342_), .Y(_2059_) );
	OAI21X1 OAI21X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_5__16_), .Y(_6343_) );
	OAI21X1 OAI21X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf3), .B(_6326__bF_buf3), .C(_6343_), .Y(_2060_) );
	OAI21X1 OAI21X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_5__17_), .Y(_6344_) );
	OAI21X1 OAI21X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf3), .B(_6326__bF_buf2), .C(_6344_), .Y(_2061_) );
	OAI21X1 OAI21X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_5__18_), .Y(_6345_) );
	OAI21X1 OAI21X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf3), .B(_6326__bF_buf1), .C(_6345_), .Y(_2062_) );
	OAI21X1 OAI21X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf12), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_5__19_), .Y(_6346_) );
	OAI21X1 OAI21X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf3), .B(_6326__bF_buf0), .C(_6346_), .Y(_2063_) );
	OAI21X1 OAI21X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf11), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_5__20_), .Y(_6347_) );
	OAI21X1 OAI21X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf3), .B(_6326__bF_buf4), .C(_6347_), .Y(_2064_) );
	OAI21X1 OAI21X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf10), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_5__21_), .Y(_6348_) );
	OAI21X1 OAI21X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf3), .B(_6326__bF_buf3), .C(_6348_), .Y(_2065_) );
	OAI21X1 OAI21X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf9), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_5__22_), .Y(_6349_) );
	OAI21X1 OAI21X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf3), .B(_6326__bF_buf2), .C(_6349_), .Y(_2066_) );
	OAI21X1 OAI21X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf8), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_5__23_), .Y(_6350_) );
	OAI21X1 OAI21X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf3), .B(_6326__bF_buf1), .C(_6350_), .Y(_2067_) );
	OAI21X1 OAI21X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf7), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_5__24_), .Y(_6351_) );
	OAI21X1 OAI21X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf3), .B(_6326__bF_buf0), .C(_6351_), .Y(_2068_) );
	OAI21X1 OAI21X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf6), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_5__25_), .Y(_6352_) );
	OAI21X1 OAI21X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf3), .B(_6326__bF_buf4), .C(_6352_), .Y(_2069_) );
	OAI21X1 OAI21X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf5), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_5__26_), .Y(_6353_) );
	OAI21X1 OAI21X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf3), .B(_6326__bF_buf3), .C(_6353_), .Y(_2070_) );
	OAI21X1 OAI21X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf4), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_5__27_), .Y(_6354_) );
	OAI21X1 OAI21X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf3), .B(_6326__bF_buf2), .C(_6354_), .Y(_2071_) );
	OAI21X1 OAI21X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf3), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_5__28_), .Y(_6355_) );
	OAI21X1 OAI21X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf3), .B(_6326__bF_buf1), .C(_6355_), .Y(_2072_) );
	OAI21X1 OAI21X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf2), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_5__29_), .Y(_6356_) );
	OAI21X1 OAI21X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf3), .B(_6326__bF_buf0), .C(_6356_), .Y(_2073_) );
	OAI21X1 OAI21X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf1), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_5__30_), .Y(_6357_) );
	OAI21X1 OAI21X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_6326__bF_buf4), .C(_6357_), .Y(_2074_) );
	OAI21X1 OAI21X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_2484__bF_buf0), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_5__31_), .Y(_6358_) );
	OAI21X1 OAI21X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf3), .B(_6326__bF_buf3), .C(_6358_), .Y(_2075_) );
	NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_6158_), .C(_2588__bF_buf3), .Y(_6359_) );
	OAI21X1 OAI21X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_6__0_), .Y(_6360_) );
	OAI21X1 OAI21X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf2), .B(_6359__bF_buf4), .C(_6360_), .Y(_2076_) );
	OAI21X1 OAI21X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_6__1_), .Y(_6361_) );
	OAI21X1 OAI21X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf2), .B(_6359__bF_buf3), .C(_6361_), .Y(_2077_) );
	OAI21X1 OAI21X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_6__2_), .Y(_6362_) );
	OAI21X1 OAI21X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf2), .B(_6359__bF_buf2), .C(_6362_), .Y(_2078_) );
	OAI21X1 OAI21X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_6__3_), .Y(_6363_) );
	OAI21X1 OAI21X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf2), .B(_6359__bF_buf1), .C(_6363_), .Y(_2079_) );
	OAI21X1 OAI21X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_6__4_), .Y(_6364_) );
	OAI21X1 OAI21X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf2), .B(_6359__bF_buf0), .C(_6364_), .Y(_2080_) );
	OAI21X1 OAI21X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_6__5_), .Y(_6365_) );
	OAI21X1 OAI21X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf2), .B(_6359__bF_buf4), .C(_6365_), .Y(_2081_) );
	OAI21X1 OAI21X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_6__6_), .Y(_6366_) );
	OAI21X1 OAI21X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf2), .B(_6359__bF_buf3), .C(_6366_), .Y(_2082_) );
	OAI21X1 OAI21X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_6__7_), .Y(_6367_) );
	OAI21X1 OAI21X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf2), .B(_6359__bF_buf2), .C(_6367_), .Y(_2083_) );
	OAI21X1 OAI21X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_6__8_), .Y(_6368_) );
	OAI21X1 OAI21X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf2), .B(_6359__bF_buf1), .C(_6368_), .Y(_2084_) );
	OAI21X1 OAI21X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_6__9_), .Y(_6369_) );
	OAI21X1 OAI21X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf2), .B(_6359__bF_buf0), .C(_6369_), .Y(_2085_) );
	OAI21X1 OAI21X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_6__10_), .Y(_6370_) );
	OAI21X1 OAI21X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf2), .B(_6359__bF_buf4), .C(_6370_), .Y(_2086_) );
	OAI21X1 OAI21X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_6__11_), .Y(_6371_) );
	OAI21X1 OAI21X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf2), .B(_6359__bF_buf3), .C(_6371_), .Y(_2087_) );
	OAI21X1 OAI21X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_6__12_), .Y(_6372_) );
	OAI21X1 OAI21X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf2), .B(_6359__bF_buf2), .C(_6372_), .Y(_2088_) );
	OAI21X1 OAI21X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_6__13_), .Y(_6373_) );
	OAI21X1 OAI21X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf2), .B(_6359__bF_buf1), .C(_6373_), .Y(_2089_) );
	OAI21X1 OAI21X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_6__14_), .Y(_6374_) );
	OAI21X1 OAI21X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf2), .B(_6359__bF_buf0), .C(_6374_), .Y(_2090_) );
	OAI21X1 OAI21X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_6__15_), .Y(_6375_) );
	OAI21X1 OAI21X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf2), .B(_6359__bF_buf4), .C(_6375_), .Y(_2091_) );
	OAI21X1 OAI21X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_6__16_), .Y(_6376_) );
	OAI21X1 OAI21X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf2), .B(_6359__bF_buf3), .C(_6376_), .Y(_2092_) );
	OAI21X1 OAI21X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_6__17_), .Y(_6377_) );
	OAI21X1 OAI21X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf2), .B(_6359__bF_buf2), .C(_6377_), .Y(_2093_) );
	OAI21X1 OAI21X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_6__18_), .Y(_6378_) );
	OAI21X1 OAI21X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf2), .B(_6359__bF_buf1), .C(_6378_), .Y(_2094_) );
	OAI21X1 OAI21X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf6), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_6__19_), .Y(_6379_) );
	OAI21X1 OAI21X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf2), .B(_6359__bF_buf0), .C(_6379_), .Y(_2095_) );
	OAI21X1 OAI21X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf5), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_6__20_), .Y(_6380_) );
	OAI21X1 OAI21X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf2), .B(_6359__bF_buf4), .C(_6380_), .Y(_2096_) );
	OAI21X1 OAI21X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf4), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_6__21_), .Y(_6381_) );
	OAI21X1 OAI21X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf2), .B(_6359__bF_buf3), .C(_6381_), .Y(_2097_) );
	OAI21X1 OAI21X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf3), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_6__22_), .Y(_6382_) );
	OAI21X1 OAI21X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf2), .B(_6359__bF_buf2), .C(_6382_), .Y(_2098_) );
	OAI21X1 OAI21X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf2), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_6__23_), .Y(_6383_) );
	OAI21X1 OAI21X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf2), .B(_6359__bF_buf1), .C(_6383_), .Y(_2099_) );
	OAI21X1 OAI21X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf1), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_6__24_), .Y(_6384_) );
	OAI21X1 OAI21X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf2), .B(_6359__bF_buf0), .C(_6384_), .Y(_2100_) );
	OAI21X1 OAI21X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf0), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_6__25_), .Y(_6385_) );
	OAI21X1 OAI21X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf2), .B(_6359__bF_buf4), .C(_6385_), .Y(_2101_) );
	OAI21X1 OAI21X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf12), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_6__26_), .Y(_6386_) );
	OAI21X1 OAI21X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf2), .B(_6359__bF_buf3), .C(_6386_), .Y(_2102_) );
	OAI21X1 OAI21X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf11), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_6__27_), .Y(_6387_) );
	OAI21X1 OAI21X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf2), .B(_6359__bF_buf2), .C(_6387_), .Y(_2103_) );
	OAI21X1 OAI21X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf10), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_6__28_), .Y(_6388_) );
	OAI21X1 OAI21X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf2), .B(_6359__bF_buf1), .C(_6388_), .Y(_2104_) );
	OAI21X1 OAI21X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf9), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_6__29_), .Y(_6389_) );
	OAI21X1 OAI21X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf2), .B(_6359__bF_buf0), .C(_6389_), .Y(_2105_) );
	OAI21X1 OAI21X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf8), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_6__30_), .Y(_6390_) );
	OAI21X1 OAI21X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_6359__bF_buf4), .C(_6390_), .Y(_2106_) );
	OAI21X1 OAI21X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_2590__bF_buf7), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_6__31_), .Y(_6391_) );
	OAI21X1 OAI21X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf2), .B(_6359__bF_buf3), .C(_6391_), .Y(_2107_) );
	NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_6158_), .C(_2623_), .Y(_6392_) );
	OAI21X1 OAI21X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_7__0_), .Y(_6393_) );
	OAI21X1 OAI21X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf1), .B(_6392__bF_buf4), .C(_6393_), .Y(_2108_) );
	OAI21X1 OAI21X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_7__1_), .Y(_6394_) );
	OAI21X1 OAI21X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf1), .B(_6392__bF_buf3), .C(_6394_), .Y(_2109_) );
	OAI21X1 OAI21X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_7__2_), .Y(_6395_) );
	OAI21X1 OAI21X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf1), .B(_6392__bF_buf2), .C(_6395_), .Y(_2110_) );
	OAI21X1 OAI21X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_7__3_), .Y(_6396_) );
	OAI21X1 OAI21X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf1), .B(_6392__bF_buf1), .C(_6396_), .Y(_2111_) );
	OAI21X1 OAI21X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_7__4_), .Y(_6397_) );
	OAI21X1 OAI21X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf1), .B(_6392__bF_buf0), .C(_6397_), .Y(_2112_) );
	OAI21X1 OAI21X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_7__5_), .Y(_6398_) );
	OAI21X1 OAI21X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf1), .B(_6392__bF_buf4), .C(_6398_), .Y(_2113_) );
	OAI21X1 OAI21X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_7__6_), .Y(_6399_) );
	OAI21X1 OAI21X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf1), .B(_6392__bF_buf3), .C(_6399_), .Y(_2114_) );
	OAI21X1 OAI21X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_7__7_), .Y(_6400_) );
	OAI21X1 OAI21X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf1), .B(_6392__bF_buf2), .C(_6400_), .Y(_2115_) );
	OAI21X1 OAI21X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_7__8_), .Y(_6401_) );
	OAI21X1 OAI21X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf1), .B(_6392__bF_buf1), .C(_6401_), .Y(_2116_) );
	OAI21X1 OAI21X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_7__9_), .Y(_6402_) );
	OAI21X1 OAI21X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf1), .B(_6392__bF_buf0), .C(_6402_), .Y(_2117_) );
	OAI21X1 OAI21X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_7__10_), .Y(_6403_) );
	OAI21X1 OAI21X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf1), .B(_6392__bF_buf4), .C(_6403_), .Y(_2118_) );
	OAI21X1 OAI21X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_7__11_), .Y(_6404_) );
	OAI21X1 OAI21X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf1), .B(_6392__bF_buf3), .C(_6404_), .Y(_2119_) );
	OAI21X1 OAI21X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_7__12_), .Y(_6405_) );
	OAI21X1 OAI21X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf1), .B(_6392__bF_buf2), .C(_6405_), .Y(_2120_) );
	OAI21X1 OAI21X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_7__13_), .Y(_6406_) );
	OAI21X1 OAI21X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf1), .B(_6392__bF_buf1), .C(_6406_), .Y(_2121_) );
	OAI21X1 OAI21X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_7__14_), .Y(_6407_) );
	OAI21X1 OAI21X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf1), .B(_6392__bF_buf0), .C(_6407_), .Y(_2122_) );
	OAI21X1 OAI21X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_7__15_), .Y(_6408_) );
	OAI21X1 OAI21X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf1), .B(_6392__bF_buf4), .C(_6408_), .Y(_2123_) );
	OAI21X1 OAI21X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_7__16_), .Y(_6409_) );
	OAI21X1 OAI21X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf1), .B(_6392__bF_buf3), .C(_6409_), .Y(_2124_) );
	OAI21X1 OAI21X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_7__17_), .Y(_6410_) );
	OAI21X1 OAI21X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf1), .B(_6392__bF_buf2), .C(_6410_), .Y(_2125_) );
	OAI21X1 OAI21X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_7__18_), .Y(_6411_) );
	OAI21X1 OAI21X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf1), .B(_6392__bF_buf1), .C(_6411_), .Y(_2126_) );
	OAI21X1 OAI21X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_7__19_), .Y(_6412_) );
	OAI21X1 OAI21X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf1), .B(_6392__bF_buf0), .C(_6412_), .Y(_2127_) );
	OAI21X1 OAI21X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_7__20_), .Y(_6413_) );
	OAI21X1 OAI21X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf1), .B(_6392__bF_buf4), .C(_6413_), .Y(_2128_) );
	OAI21X1 OAI21X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6293__bF_buf3), .C(csr_gpr_iu_gpr_7__21_), .Y(_6414_) );
	OAI21X1 OAI21X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf1), .B(_6392__bF_buf3), .C(_6414_), .Y(_2129_) );
	OAI21X1 OAI21X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6293__bF_buf2), .C(csr_gpr_iu_gpr_7__22_), .Y(_6415_) );
	OAI21X1 OAI21X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf1), .B(_6392__bF_buf2), .C(_6415_), .Y(_2130_) );
	OAI21X1 OAI21X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6293__bF_buf1), .C(csr_gpr_iu_gpr_7__23_), .Y(_6416_) );
	OAI21X1 OAI21X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf1), .B(_6392__bF_buf1), .C(_6416_), .Y(_2131_) );
	OAI21X1 OAI21X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6293__bF_buf0), .C(csr_gpr_iu_gpr_7__24_), .Y(_6417_) );
	OAI21X1 OAI21X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf1), .B(_6392__bF_buf0), .C(_6417_), .Y(_2132_) );
	OAI21X1 OAI21X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6293__bF_buf10), .C(csr_gpr_iu_gpr_7__25_), .Y(_6418_) );
	OAI21X1 OAI21X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf1), .B(_6392__bF_buf4), .C(_6418_), .Y(_2133_) );
	OAI21X1 OAI21X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6293__bF_buf9), .C(csr_gpr_iu_gpr_7__26_), .Y(_6419_) );
	OAI21X1 OAI21X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf1), .B(_6392__bF_buf3), .C(_6419_), .Y(_2134_) );
	OAI21X1 OAI21X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6293__bF_buf8), .C(csr_gpr_iu_gpr_7__27_), .Y(_6420_) );
	OAI21X1 OAI21X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf1), .B(_6392__bF_buf2), .C(_6420_), .Y(_2135_) );
	OAI21X1 OAI21X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6293__bF_buf7), .C(csr_gpr_iu_gpr_7__28_), .Y(_6421_) );
	OAI21X1 OAI21X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf1), .B(_6392__bF_buf1), .C(_6421_), .Y(_2136_) );
	OAI21X1 OAI21X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6293__bF_buf6), .C(csr_gpr_iu_gpr_7__29_), .Y(_6422_) );
	OAI21X1 OAI21X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf1), .B(_6392__bF_buf0), .C(_6422_), .Y(_2137_) );
	OAI21X1 OAI21X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6293__bF_buf5), .C(csr_gpr_iu_gpr_7__30_), .Y(_6423_) );
	OAI21X1 OAI21X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_6392__bF_buf4), .C(_6423_), .Y(_2138_) );
	OAI21X1 OAI21X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6293__bF_buf4), .C(csr_gpr_iu_gpr_7__31_), .Y(_6424_) );
	OAI21X1 OAI21X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf1), .B(_6392__bF_buf3), .C(_6424_), .Y(_2139_) );
	NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2694__bF_buf3), .C(_6024_), .Y(_6425_) );
	NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2551_), .C(_2476_), .Y(_6426_) );
	OAI21X1 OAI21X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2696__bF_buf12), .C(csr_gpr_iu_gpr_8__0_), .Y(_6427_) );
	OAI21X1 OAI21X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf0), .B(_6425__bF_buf4), .C(_6427_), .Y(_2140_) );
	OAI21X1 OAI21X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2696__bF_buf11), .C(csr_gpr_iu_gpr_8__1_), .Y(_6428_) );
	OAI21X1 OAI21X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf0), .B(_6425__bF_buf3), .C(_6428_), .Y(_2141_) );
	OAI21X1 OAI21X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2696__bF_buf10), .C(csr_gpr_iu_gpr_8__2_), .Y(_6429_) );
	OAI21X1 OAI21X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf0), .B(_6425__bF_buf2), .C(_6429_), .Y(_2142_) );
	OAI21X1 OAI21X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2696__bF_buf9), .C(csr_gpr_iu_gpr_8__3_), .Y(_6430_) );
	OAI21X1 OAI21X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf0), .B(_6425__bF_buf1), .C(_6430_), .Y(_2143_) );
	OAI21X1 OAI21X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2696__bF_buf8), .C(csr_gpr_iu_gpr_8__4_), .Y(_6431_) );
	OAI21X1 OAI21X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf0), .B(_6425__bF_buf0), .C(_6431_), .Y(_2144_) );
	OAI21X1 OAI21X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2696__bF_buf7), .C(csr_gpr_iu_gpr_8__5_), .Y(_6432_) );
	OAI21X1 OAI21X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf0), .B(_6425__bF_buf4), .C(_6432_), .Y(_2145_) );
	OAI21X1 OAI21X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2696__bF_buf6), .C(csr_gpr_iu_gpr_8__6_), .Y(_6433_) );
	OAI21X1 OAI21X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf0), .B(_6425__bF_buf3), .C(_6433_), .Y(_2146_) );
	OAI21X1 OAI21X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2696__bF_buf5), .C(csr_gpr_iu_gpr_8__7_), .Y(_6434_) );
	OAI21X1 OAI21X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf0), .B(_6425__bF_buf2), .C(_6434_), .Y(_2147_) );
	OAI21X1 OAI21X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2696__bF_buf4), .C(csr_gpr_iu_gpr_8__8_), .Y(_6435_) );
	OAI21X1 OAI21X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf0), .B(_6425__bF_buf1), .C(_6435_), .Y(_2148_) );
	OAI21X1 OAI21X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2696__bF_buf3), .C(csr_gpr_iu_gpr_8__9_), .Y(_6436_) );
	OAI21X1 OAI21X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf0), .B(_6425__bF_buf0), .C(_6436_), .Y(_2149_) );
	OAI21X1 OAI21X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2696__bF_buf2), .C(csr_gpr_iu_gpr_8__10_), .Y(_6437_) );
	OAI21X1 OAI21X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf0), .B(_6425__bF_buf4), .C(_6437_), .Y(_2150_) );
	OAI21X1 OAI21X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2696__bF_buf1), .C(csr_gpr_iu_gpr_8__11_), .Y(_6438_) );
	OAI21X1 OAI21X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf0), .B(_6425__bF_buf3), .C(_6438_), .Y(_2151_) );
	OAI21X1 OAI21X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2696__bF_buf0), .C(csr_gpr_iu_gpr_8__12_), .Y(_6439_) );
	OAI21X1 OAI21X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf0), .B(_6425__bF_buf2), .C(_6439_), .Y(_2152_) );
	OAI21X1 OAI21X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2696__bF_buf12), .C(csr_gpr_iu_gpr_8__13_), .Y(_6440_) );
	OAI21X1 OAI21X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf0), .B(_6425__bF_buf1), .C(_6440_), .Y(_2153_) );
	OAI21X1 OAI21X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2696__bF_buf11), .C(csr_gpr_iu_gpr_8__14_), .Y(_6441_) );
	OAI21X1 OAI21X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf0), .B(_6425__bF_buf0), .C(_6441_), .Y(_2154_) );
	OAI21X1 OAI21X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2696__bF_buf10), .C(csr_gpr_iu_gpr_8__15_), .Y(_6442_) );
	OAI21X1 OAI21X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf0), .B(_6425__bF_buf4), .C(_6442_), .Y(_2155_) );
	OAI21X1 OAI21X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2696__bF_buf9), .C(csr_gpr_iu_gpr_8__16_), .Y(_6443_) );
	OAI21X1 OAI21X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf0), .B(_6425__bF_buf3), .C(_6443_), .Y(_2156_) );
	OAI21X1 OAI21X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2696__bF_buf8), .C(csr_gpr_iu_gpr_8__17_), .Y(_6444_) );
	OAI21X1 OAI21X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf0), .B(_6425__bF_buf2), .C(_6444_), .Y(_2157_) );
	OAI21X1 OAI21X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2696__bF_buf7), .C(csr_gpr_iu_gpr_8__18_), .Y(_6445_) );
	OAI21X1 OAI21X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf0), .B(_6425__bF_buf1), .C(_6445_), .Y(_2158_) );
	OAI21X1 OAI21X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2696__bF_buf6), .C(csr_gpr_iu_gpr_8__19_), .Y(_6446_) );
	OAI21X1 OAI21X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf0), .B(_6425__bF_buf0), .C(_6446_), .Y(_2159_) );
	OAI21X1 OAI21X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2696__bF_buf5), .C(csr_gpr_iu_gpr_8__20_), .Y(_6447_) );
	OAI21X1 OAI21X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf0), .B(_6425__bF_buf4), .C(_6447_), .Y(_2160_) );
	OAI21X1 OAI21X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2696__bF_buf4), .C(csr_gpr_iu_gpr_8__21_), .Y(_6448_) );
	OAI21X1 OAI21X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf0), .B(_6425__bF_buf3), .C(_6448_), .Y(_2161_) );
	OAI21X1 OAI21X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2696__bF_buf3), .C(csr_gpr_iu_gpr_8__22_), .Y(_6449_) );
	OAI21X1 OAI21X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf0), .B(_6425__bF_buf2), .C(_6449_), .Y(_2162_) );
	OAI21X1 OAI21X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2696__bF_buf2), .C(csr_gpr_iu_gpr_8__23_), .Y(_6450_) );
	OAI21X1 OAI21X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf0), .B(_6425__bF_buf1), .C(_6450_), .Y(_2163_) );
	OAI21X1 OAI21X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2696__bF_buf1), .C(csr_gpr_iu_gpr_8__24_), .Y(_6451_) );
	OAI21X1 OAI21X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf0), .B(_6425__bF_buf0), .C(_6451_), .Y(_2164_) );
	OAI21X1 OAI21X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2696__bF_buf0), .C(csr_gpr_iu_gpr_8__25_), .Y(_6452_) );
	OAI21X1 OAI21X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf0), .B(_6425__bF_buf4), .C(_6452_), .Y(_2165_) );
	OAI21X1 OAI21X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2696__bF_buf12), .C(csr_gpr_iu_gpr_8__26_), .Y(_6453_) );
	OAI21X1 OAI21X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf0), .B(_6425__bF_buf3), .C(_6453_), .Y(_2166_) );
	OAI21X1 OAI21X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2696__bF_buf11), .C(csr_gpr_iu_gpr_8__27_), .Y(_6454_) );
	OAI21X1 OAI21X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf0), .B(_6425__bF_buf2), .C(_6454_), .Y(_2167_) );
	OAI21X1 OAI21X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2696__bF_buf10), .C(csr_gpr_iu_gpr_8__28_), .Y(_6455_) );
	OAI21X1 OAI21X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf0), .B(_6425__bF_buf1), .C(_6455_), .Y(_2168_) );
	OAI21X1 OAI21X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2696__bF_buf9), .C(csr_gpr_iu_gpr_8__29_), .Y(_6456_) );
	OAI21X1 OAI21X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf0), .B(_6425__bF_buf0), .C(_6456_), .Y(_2169_) );
	OAI21X1 OAI21X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2696__bF_buf8), .C(csr_gpr_iu_gpr_8__30_), .Y(_6457_) );
	OAI21X1 OAI21X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_6425__bF_buf4), .C(_6457_), .Y(_2170_) );
	OAI21X1 OAI21X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2696__bF_buf7), .C(csr_gpr_iu_gpr_8__31_), .Y(_6458_) );
	OAI21X1 OAI21X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf0), .B(_6425__bF_buf3), .C(_6458_), .Y(_2171_) );
	NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2694__bF_buf2), .C(_6024_), .Y(_6459_) );
	OAI21X1 OAI21X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2696__bF_buf6), .C(csr_gpr_iu_gpr_12__0_), .Y(_6460_) );
	OAI21X1 OAI21X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf4), .B(_6459__bF_buf4), .C(_6460_), .Y(_2172_) );
	OAI21X1 OAI21X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2696__bF_buf5), .C(csr_gpr_iu_gpr_12__1_), .Y(_6461_) );
	OAI21X1 OAI21X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf4), .B(_6459__bF_buf3), .C(_6461_), .Y(_2173_) );
	OAI21X1 OAI21X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2696__bF_buf4), .C(csr_gpr_iu_gpr_12__2_), .Y(_6462_) );
	OAI21X1 OAI21X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf4), .B(_6459__bF_buf2), .C(_6462_), .Y(_2174_) );
	OAI21X1 OAI21X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2696__bF_buf3), .C(csr_gpr_iu_gpr_12__3_), .Y(_6463_) );
	OAI21X1 OAI21X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf4), .B(_6459__bF_buf1), .C(_6463_), .Y(_2175_) );
	OAI21X1 OAI21X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2696__bF_buf2), .C(csr_gpr_iu_gpr_12__4_), .Y(_6464_) );
	OAI21X1 OAI21X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf4), .B(_6459__bF_buf0), .C(_6464_), .Y(_2176_) );
	OAI21X1 OAI21X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2696__bF_buf1), .C(csr_gpr_iu_gpr_12__5_), .Y(_6465_) );
	OAI21X1 OAI21X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf4), .B(_6459__bF_buf4), .C(_6465_), .Y(_2177_) );
	OAI21X1 OAI21X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2696__bF_buf0), .C(csr_gpr_iu_gpr_12__6_), .Y(_6466_) );
	OAI21X1 OAI21X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf4), .B(_6459__bF_buf3), .C(_6466_), .Y(_2178_) );
	OAI21X1 OAI21X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2696__bF_buf12), .C(csr_gpr_iu_gpr_12__7_), .Y(_6467_) );
	OAI21X1 OAI21X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf4), .B(_6459__bF_buf2), .C(_6467_), .Y(_2179_) );
	OAI21X1 OAI21X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2696__bF_buf11), .C(csr_gpr_iu_gpr_12__8_), .Y(_6468_) );
	OAI21X1 OAI21X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf4), .B(_6459__bF_buf1), .C(_6468_), .Y(_2180_) );
	OAI21X1 OAI21X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2696__bF_buf10), .C(csr_gpr_iu_gpr_12__9_), .Y(_6469_) );
	OAI21X1 OAI21X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf4), .B(_6459__bF_buf0), .C(_6469_), .Y(_2181_) );
	OAI21X1 OAI21X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2696__bF_buf9), .C(csr_gpr_iu_gpr_12__10_), .Y(_6470_) );
	OAI21X1 OAI21X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf4), .B(_6459__bF_buf4), .C(_6470_), .Y(_2182_) );
	OAI21X1 OAI21X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2696__bF_buf8), .C(csr_gpr_iu_gpr_12__11_), .Y(_6471_) );
	OAI21X1 OAI21X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf4), .B(_6459__bF_buf3), .C(_6471_), .Y(_2183_) );
	OAI21X1 OAI21X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2696__bF_buf7), .C(csr_gpr_iu_gpr_12__12_), .Y(_6472_) );
	OAI21X1 OAI21X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf4), .B(_6459__bF_buf2), .C(_6472_), .Y(_2184_) );
	OAI21X1 OAI21X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2696__bF_buf6), .C(csr_gpr_iu_gpr_12__13_), .Y(_6473_) );
	OAI21X1 OAI21X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf4), .B(_6459__bF_buf1), .C(_6473_), .Y(_2185_) );
	OAI21X1 OAI21X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2696__bF_buf5), .C(csr_gpr_iu_gpr_12__14_), .Y(_6474_) );
	OAI21X1 OAI21X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf4), .B(_6459__bF_buf0), .C(_6474_), .Y(_2186_) );
	OAI21X1 OAI21X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2696__bF_buf4), .C(csr_gpr_iu_gpr_12__15_), .Y(_6475_) );
	OAI21X1 OAI21X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf4), .B(_6459__bF_buf4), .C(_6475_), .Y(_2187_) );
	OAI21X1 OAI21X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2696__bF_buf3), .C(csr_gpr_iu_gpr_12__16_), .Y(_6476_) );
	OAI21X1 OAI21X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf4), .B(_6459__bF_buf3), .C(_6476_), .Y(_2188_) );
	OAI21X1 OAI21X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2696__bF_buf2), .C(csr_gpr_iu_gpr_12__17_), .Y(_6477_) );
	OAI21X1 OAI21X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf4), .B(_6459__bF_buf2), .C(_6477_), .Y(_2189_) );
	OAI21X1 OAI21X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2696__bF_buf1), .C(csr_gpr_iu_gpr_12__18_), .Y(_6478_) );
	OAI21X1 OAI21X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf4), .B(_6459__bF_buf1), .C(_6478_), .Y(_2190_) );
	OAI21X1 OAI21X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2696__bF_buf0), .C(csr_gpr_iu_gpr_12__19_), .Y(_6479_) );
	OAI21X1 OAI21X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf4), .B(_6459__bF_buf0), .C(_6479_), .Y(_2191_) );
	OAI21X1 OAI21X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2696__bF_buf12), .C(csr_gpr_iu_gpr_12__20_), .Y(_6480_) );
	OAI21X1 OAI21X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf4), .B(_6459__bF_buf4), .C(_6480_), .Y(_2192_) );
	OAI21X1 OAI21X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2696__bF_buf11), .C(csr_gpr_iu_gpr_12__21_), .Y(_6481_) );
	OAI21X1 OAI21X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf4), .B(_6459__bF_buf3), .C(_6481_), .Y(_2193_) );
	OAI21X1 OAI21X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2696__bF_buf10), .C(csr_gpr_iu_gpr_12__22_), .Y(_6482_) );
	OAI21X1 OAI21X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf4), .B(_6459__bF_buf2), .C(_6482_), .Y(_2194_) );
	OAI21X1 OAI21X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2696__bF_buf9), .C(csr_gpr_iu_gpr_12__23_), .Y(_6483_) );
	OAI21X1 OAI21X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf4), .B(_6459__bF_buf1), .C(_6483_), .Y(_2195_) );
	OAI21X1 OAI21X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2696__bF_buf8), .C(csr_gpr_iu_gpr_12__24_), .Y(_6484_) );
	OAI21X1 OAI21X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf4), .B(_6459__bF_buf0), .C(_6484_), .Y(_2196_) );
	OAI21X1 OAI21X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2696__bF_buf7), .C(csr_gpr_iu_gpr_12__25_), .Y(_6485_) );
	OAI21X1 OAI21X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf4), .B(_6459__bF_buf4), .C(_6485_), .Y(_2197_) );
	OAI21X1 OAI21X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2696__bF_buf6), .C(csr_gpr_iu_gpr_12__26_), .Y(_6486_) );
	OAI21X1 OAI21X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf4), .B(_6459__bF_buf3), .C(_6486_), .Y(_2198_) );
	OAI21X1 OAI21X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2696__bF_buf5), .C(csr_gpr_iu_gpr_12__27_), .Y(_6487_) );
	OAI21X1 OAI21X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf4), .B(_6459__bF_buf2), .C(_6487_), .Y(_2199_) );
	OAI21X1 OAI21X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2696__bF_buf4), .C(csr_gpr_iu_gpr_12__28_), .Y(_6488_) );
	OAI21X1 OAI21X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf4), .B(_6459__bF_buf1), .C(_6488_), .Y(_2200_) );
	OAI21X1 OAI21X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2696__bF_buf3), .C(csr_gpr_iu_gpr_12__29_), .Y(_6489_) );
	OAI21X1 OAI21X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf4), .B(_6459__bF_buf0), .C(_6489_), .Y(_2201_) );
	OAI21X1 OAI21X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2696__bF_buf2), .C(csr_gpr_iu_gpr_12__30_), .Y(_6490_) );
	OAI21X1 OAI21X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_6459__bF_buf4), .C(_6490_), .Y(_2202_) );
	OAI21X1 OAI21X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2696__bF_buf1), .C(csr_gpr_iu_gpr_12__31_), .Y(_6491_) );
	OAI21X1 OAI21X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf4), .B(_6459__bF_buf3), .C(_6491_), .Y(_2203_) );
	NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2473__bF_buf3), .C(_6024_), .Y(_6492_) );
	OAI21X1 OAI21X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2484__bF_buf12), .C(csr_gpr_iu_gpr_13__0_), .Y(_6493_) );
	OAI21X1 OAI21X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf3), .B(_6492__bF_buf4), .C(_6493_), .Y(_2204_) );
	OAI21X1 OAI21X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2484__bF_buf11), .C(csr_gpr_iu_gpr_13__1_), .Y(_6494_) );
	OAI21X1 OAI21X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf3), .B(_6492__bF_buf3), .C(_6494_), .Y(_2205_) );
	OAI21X1 OAI21X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2484__bF_buf10), .C(csr_gpr_iu_gpr_13__2_), .Y(_6495_) );
	OAI21X1 OAI21X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf3), .B(_6492__bF_buf2), .C(_6495_), .Y(_2206_) );
	OAI21X1 OAI21X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2484__bF_buf9), .C(csr_gpr_iu_gpr_13__3_), .Y(_6496_) );
	OAI21X1 OAI21X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf3), .B(_6492__bF_buf1), .C(_6496_), .Y(_2207_) );
	OAI21X1 OAI21X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2484__bF_buf8), .C(csr_gpr_iu_gpr_13__4_), .Y(_6497_) );
	OAI21X1 OAI21X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf3), .B(_6492__bF_buf0), .C(_6497_), .Y(_2208_) );
	OAI21X1 OAI21X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2484__bF_buf7), .C(csr_gpr_iu_gpr_13__5_), .Y(_6498_) );
	OAI21X1 OAI21X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf3), .B(_6492__bF_buf4), .C(_6498_), .Y(_2209_) );
	OAI21X1 OAI21X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2484__bF_buf6), .C(csr_gpr_iu_gpr_13__6_), .Y(_6499_) );
	OAI21X1 OAI21X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf3), .B(_6492__bF_buf3), .C(_6499_), .Y(_2210_) );
	OAI21X1 OAI21X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2484__bF_buf5), .C(csr_gpr_iu_gpr_13__7_), .Y(_6500_) );
	OAI21X1 OAI21X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf3), .B(_6492__bF_buf2), .C(_6500_), .Y(_2211_) );
	OAI21X1 OAI21X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2484__bF_buf4), .C(csr_gpr_iu_gpr_13__8_), .Y(_6501_) );
	OAI21X1 OAI21X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf3), .B(_6492__bF_buf1), .C(_6501_), .Y(_2212_) );
	OAI21X1 OAI21X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2484__bF_buf3), .C(csr_gpr_iu_gpr_13__9_), .Y(_6502_) );
	OAI21X1 OAI21X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf3), .B(_6492__bF_buf0), .C(_6502_), .Y(_2213_) );
	OAI21X1 OAI21X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2484__bF_buf2), .C(csr_gpr_iu_gpr_13__10_), .Y(_6503_) );
	OAI21X1 OAI21X1_2921 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf3), .B(_6492__bF_buf4), .C(_6503_), .Y(_2214_) );
	OAI21X1 OAI21X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2484__bF_buf1), .C(csr_gpr_iu_gpr_13__11_), .Y(_6504_) );
	OAI21X1 OAI21X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf3), .B(_6492__bF_buf3), .C(_6504_), .Y(_2215_) );
	OAI21X1 OAI21X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2484__bF_buf0), .C(csr_gpr_iu_gpr_13__12_), .Y(_6505_) );
	OAI21X1 OAI21X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf3), .B(_6492__bF_buf2), .C(_6505_), .Y(_2216_) );
	OAI21X1 OAI21X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2484__bF_buf12), .C(csr_gpr_iu_gpr_13__13_), .Y(_6506_) );
	OAI21X1 OAI21X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf3), .B(_6492__bF_buf1), .C(_6506_), .Y(_2217_) );
	OAI21X1 OAI21X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2484__bF_buf11), .C(csr_gpr_iu_gpr_13__14_), .Y(_6507_) );
	OAI21X1 OAI21X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf3), .B(_6492__bF_buf0), .C(_6507_), .Y(_2218_) );
	OAI21X1 OAI21X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2484__bF_buf10), .C(csr_gpr_iu_gpr_13__15_), .Y(_6508_) );
	OAI21X1 OAI21X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf3), .B(_6492__bF_buf4), .C(_6508_), .Y(_2219_) );
	OAI21X1 OAI21X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2484__bF_buf9), .C(csr_gpr_iu_gpr_13__16_), .Y(_6509_) );
	OAI21X1 OAI21X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf3), .B(_6492__bF_buf3), .C(_6509_), .Y(_2220_) );
	OAI21X1 OAI21X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2484__bF_buf8), .C(csr_gpr_iu_gpr_13__17_), .Y(_6510_) );
	OAI21X1 OAI21X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf3), .B(_6492__bF_buf2), .C(_6510_), .Y(_2221_) );
	OAI21X1 OAI21X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2484__bF_buf7), .C(csr_gpr_iu_gpr_13__18_), .Y(_6511_) );
	OAI21X1 OAI21X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf3), .B(_6492__bF_buf1), .C(_6511_), .Y(_2222_) );
	OAI21X1 OAI21X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2484__bF_buf6), .C(csr_gpr_iu_gpr_13__19_), .Y(_6512_) );
	OAI21X1 OAI21X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf3), .B(_6492__bF_buf0), .C(_6512_), .Y(_2223_) );
	OAI21X1 OAI21X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2484__bF_buf5), .C(csr_gpr_iu_gpr_13__20_), .Y(_6513_) );
	OAI21X1 OAI21X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf3), .B(_6492__bF_buf4), .C(_6513_), .Y(_2224_) );
	OAI21X1 OAI21X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf2), .B(_2484__bF_buf4), .C(csr_gpr_iu_gpr_13__21_), .Y(_6514_) );
	OAI21X1 OAI21X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf3), .B(_6492__bF_buf3), .C(_6514_), .Y(_2225_) );
	OAI21X1 OAI21X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf1), .B(_2484__bF_buf3), .C(csr_gpr_iu_gpr_13__22_), .Y(_6515_) );
	OAI21X1 OAI21X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf3), .B(_6492__bF_buf2), .C(_6515_), .Y(_2226_) );
	OAI21X1 OAI21X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf0), .B(_2484__bF_buf2), .C(csr_gpr_iu_gpr_13__23_), .Y(_6516_) );
	OAI21X1 OAI21X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf3), .B(_6492__bF_buf1), .C(_6516_), .Y(_2227_) );
	OAI21X1 OAI21X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf10), .B(_2484__bF_buf1), .C(csr_gpr_iu_gpr_13__24_), .Y(_6517_) );
	OAI21X1 OAI21X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf3), .B(_6492__bF_buf0), .C(_6517_), .Y(_2228_) );
	OAI21X1 OAI21X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf9), .B(_2484__bF_buf0), .C(csr_gpr_iu_gpr_13__25_), .Y(_6518_) );
	OAI21X1 OAI21X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf3), .B(_6492__bF_buf4), .C(_6518_), .Y(_2229_) );
	OAI21X1 OAI21X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf8), .B(_2484__bF_buf12), .C(csr_gpr_iu_gpr_13__26_), .Y(_6519_) );
	OAI21X1 OAI21X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf3), .B(_6492__bF_buf3), .C(_6519_), .Y(_2230_) );
	OAI21X1 OAI21X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf7), .B(_2484__bF_buf11), .C(csr_gpr_iu_gpr_13__27_), .Y(_6520_) );
	OAI21X1 OAI21X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf3), .B(_6492__bF_buf2), .C(_6520_), .Y(_2231_) );
	OAI21X1 OAI21X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf6), .B(_2484__bF_buf10), .C(csr_gpr_iu_gpr_13__28_), .Y(_6521_) );
	OAI21X1 OAI21X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf3), .B(_6492__bF_buf1), .C(_6521_), .Y(_2232_) );
	OAI21X1 OAI21X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf5), .B(_2484__bF_buf9), .C(csr_gpr_iu_gpr_13__29_), .Y(_6522_) );
	OAI21X1 OAI21X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf3), .B(_6492__bF_buf0), .C(_6522_), .Y(_2233_) );
	OAI21X1 OAI21X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf4), .B(_2484__bF_buf8), .C(csr_gpr_iu_gpr_13__30_), .Y(_6523_) );
	OAI21X1 OAI21X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_6492__bF_buf4), .C(_6523_), .Y(_2234_) );
	OAI21X1 OAI21X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_6026__bF_buf3), .B(_2484__bF_buf7), .C(csr_gpr_iu_gpr_13__31_), .Y(_6524_) );
	OAI21X1 OAI21X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf3), .B(_6492__bF_buf3), .C(_6524_), .Y(_2235_) );
	NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2473__bF_buf2), .C(_6024_), .Y(_6525_) );
	OAI21X1 OAI21X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2484__bF_buf6), .C(csr_gpr_iu_gpr_9__0_), .Y(_6526_) );
	OAI21X1 OAI21X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf2), .B(_6525__bF_buf4), .C(_6526_), .Y(_2236_) );
	OAI21X1 OAI21X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2484__bF_buf5), .C(csr_gpr_iu_gpr_9__1_), .Y(_6527_) );
	OAI21X1 OAI21X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf2), .B(_6525__bF_buf3), .C(_6527_), .Y(_2237_) );
	OAI21X1 OAI21X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2484__bF_buf4), .C(csr_gpr_iu_gpr_9__2_), .Y(_6528_) );
	OAI21X1 OAI21X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf2), .B(_6525__bF_buf2), .C(_6528_), .Y(_2238_) );
	OAI21X1 OAI21X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2484__bF_buf3), .C(csr_gpr_iu_gpr_9__3_), .Y(_6529_) );
	OAI21X1 OAI21X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf2), .B(_6525__bF_buf1), .C(_6529_), .Y(_2239_) );
	OAI21X1 OAI21X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2484__bF_buf2), .C(csr_gpr_iu_gpr_9__4_), .Y(_6530_) );
	OAI21X1 OAI21X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf2), .B(_6525__bF_buf0), .C(_6530_), .Y(_2240_) );
	OAI21X1 OAI21X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2484__bF_buf1), .C(csr_gpr_iu_gpr_9__5_), .Y(_6531_) );
	OAI21X1 OAI21X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf2), .B(_6525__bF_buf4), .C(_6531_), .Y(_2241_) );
	OAI21X1 OAI21X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2484__bF_buf0), .C(csr_gpr_iu_gpr_9__6_), .Y(_6532_) );
	OAI21X1 OAI21X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf2), .B(_6525__bF_buf3), .C(_6532_), .Y(_2242_) );
	OAI21X1 OAI21X1_2978 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2484__bF_buf12), .C(csr_gpr_iu_gpr_9__7_), .Y(_6533_) );
	OAI21X1 OAI21X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf2), .B(_6525__bF_buf2), .C(_6533_), .Y(_2243_) );
	OAI21X1 OAI21X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2484__bF_buf11), .C(csr_gpr_iu_gpr_9__8_), .Y(_6534_) );
	OAI21X1 OAI21X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf2), .B(_6525__bF_buf1), .C(_6534_), .Y(_2244_) );
	OAI21X1 OAI21X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2484__bF_buf10), .C(csr_gpr_iu_gpr_9__9_), .Y(_6535_) );
	OAI21X1 OAI21X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf2), .B(_6525__bF_buf0), .C(_6535_), .Y(_2245_) );
	OAI21X1 OAI21X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2484__bF_buf9), .C(csr_gpr_iu_gpr_9__10_), .Y(_6536_) );
	OAI21X1 OAI21X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf2), .B(_6525__bF_buf4), .C(_6536_), .Y(_2246_) );
	OAI21X1 OAI21X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2484__bF_buf8), .C(csr_gpr_iu_gpr_9__11_), .Y(_6537_) );
	OAI21X1 OAI21X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf2), .B(_6525__bF_buf3), .C(_6537_), .Y(_2247_) );
	OAI21X1 OAI21X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2484__bF_buf7), .C(csr_gpr_iu_gpr_9__12_), .Y(_6538_) );
	OAI21X1 OAI21X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf2), .B(_6525__bF_buf2), .C(_6538_), .Y(_2248_) );
	OAI21X1 OAI21X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2484__bF_buf6), .C(csr_gpr_iu_gpr_9__13_), .Y(_6539_) );
	OAI21X1 OAI21X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf2), .B(_6525__bF_buf1), .C(_6539_), .Y(_2249_) );
	OAI21X1 OAI21X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2484__bF_buf5), .C(csr_gpr_iu_gpr_9__14_), .Y(_6540_) );
	OAI21X1 OAI21X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf2), .B(_6525__bF_buf0), .C(_6540_), .Y(_2250_) );
	OAI21X1 OAI21X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2484__bF_buf4), .C(csr_gpr_iu_gpr_9__15_), .Y(_6541_) );
	OAI21X1 OAI21X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf2), .B(_6525__bF_buf4), .C(_6541_), .Y(_2251_) );
	OAI21X1 OAI21X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2484__bF_buf3), .C(csr_gpr_iu_gpr_9__16_), .Y(_6542_) );
	OAI21X1 OAI21X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf2), .B(_6525__bF_buf3), .C(_6542_), .Y(_2252_) );
	OAI21X1 OAI21X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2484__bF_buf2), .C(csr_gpr_iu_gpr_9__17_), .Y(_6543_) );
	OAI21X1 OAI21X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf2), .B(_6525__bF_buf2), .C(_6543_), .Y(_2253_) );
	OAI21X1 OAI21X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2484__bF_buf1), .C(csr_gpr_iu_gpr_9__18_), .Y(_6544_) );
	OAI21X1 OAI21X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf2), .B(_6525__bF_buf1), .C(_6544_), .Y(_2254_) );
	OAI21X1 OAI21X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2484__bF_buf0), .C(csr_gpr_iu_gpr_9__19_), .Y(_6545_) );
	OAI21X1 OAI21X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf2), .B(_6525__bF_buf0), .C(_6545_), .Y(_2255_) );
	OAI21X1 OAI21X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2484__bF_buf12), .C(csr_gpr_iu_gpr_9__20_), .Y(_6546_) );
	OAI21X1 OAI21X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf2), .B(_6525__bF_buf4), .C(_6546_), .Y(_2256_) );
	OAI21X1 OAI21X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2484__bF_buf11), .C(csr_gpr_iu_gpr_9__21_), .Y(_6547_) );
	OAI21X1 OAI21X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf2), .B(_6525__bF_buf3), .C(_6547_), .Y(_2257_) );
	OAI21X1 OAI21X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2484__bF_buf10), .C(csr_gpr_iu_gpr_9__22_), .Y(_6548_) );
	OAI21X1 OAI21X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf2), .B(_6525__bF_buf2), .C(_6548_), .Y(_2258_) );
	OAI21X1 OAI21X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2484__bF_buf9), .C(csr_gpr_iu_gpr_9__23_), .Y(_6549_) );
	OAI21X1 OAI21X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf2), .B(_6525__bF_buf1), .C(_6549_), .Y(_2259_) );
	OAI21X1 OAI21X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2484__bF_buf8), .C(csr_gpr_iu_gpr_9__24_), .Y(_6550_) );
	OAI21X1 OAI21X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf2), .B(_6525__bF_buf0), .C(_6550_), .Y(_2260_) );
	OAI21X1 OAI21X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2484__bF_buf7), .C(csr_gpr_iu_gpr_9__25_), .Y(_6551_) );
	OAI21X1 OAI21X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf2), .B(_6525__bF_buf4), .C(_6551_), .Y(_2261_) );
	OAI21X1 OAI21X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2484__bF_buf6), .C(csr_gpr_iu_gpr_9__26_), .Y(_6552_) );
	OAI21X1 OAI21X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf2), .B(_6525__bF_buf3), .C(_6552_), .Y(_2262_) );
	OAI21X1 OAI21X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2484__bF_buf5), .C(csr_gpr_iu_gpr_9__27_), .Y(_6553_) );
	OAI21X1 OAI21X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf2), .B(_6525__bF_buf2), .C(_6553_), .Y(_2263_) );
	OAI21X1 OAI21X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2484__bF_buf4), .C(csr_gpr_iu_gpr_9__28_), .Y(_6554_) );
	OAI21X1 OAI21X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf2), .B(_6525__bF_buf1), .C(_6554_), .Y(_2264_) );
	OAI21X1 OAI21X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2484__bF_buf3), .C(csr_gpr_iu_gpr_9__29_), .Y(_6555_) );
	OAI21X1 OAI21X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf2), .B(_6525__bF_buf0), .C(_6555_), .Y(_2265_) );
	OAI21X1 OAI21X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2484__bF_buf2), .C(csr_gpr_iu_gpr_9__30_), .Y(_6556_) );
	OAI21X1 OAI21X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_6525__bF_buf4), .C(_6556_), .Y(_2266_) );
	OAI21X1 OAI21X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2484__bF_buf1), .C(csr_gpr_iu_gpr_9__31_), .Y(_6557_) );
	OAI21X1 OAI21X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf2), .B(_6525__bF_buf3), .C(_6557_), .Y(_2267_) );
	NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2588__bF_buf2), .C(_6024_), .Y(_6558_) );
	OAI21X1 OAI21X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_10__0_), .Y(_6559_) );
	OAI21X1 OAI21X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf1), .B(_6558__bF_buf4), .C(_6559_), .Y(_2268_) );
	OAI21X1 OAI21X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2590__bF_buf5), .C(csr_gpr_iu_gpr_10__1_), .Y(_6560_) );
	OAI21X1 OAI21X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf1), .B(_6558__bF_buf3), .C(_6560_), .Y(_2269_) );
	OAI21X1 OAI21X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2590__bF_buf4), .C(csr_gpr_iu_gpr_10__2_), .Y(_6561_) );
	OAI21X1 OAI21X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf1), .B(_6558__bF_buf2), .C(_6561_), .Y(_2270_) );
	OAI21X1 OAI21X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2590__bF_buf3), .C(csr_gpr_iu_gpr_10__3_), .Y(_6562_) );
	OAI21X1 OAI21X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf1), .B(_6558__bF_buf1), .C(_6562_), .Y(_2271_) );
	OAI21X1 OAI21X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2590__bF_buf2), .C(csr_gpr_iu_gpr_10__4_), .Y(_6563_) );
	OAI21X1 OAI21X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf1), .B(_6558__bF_buf0), .C(_6563_), .Y(_2272_) );
	OAI21X1 OAI21X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2590__bF_buf1), .C(csr_gpr_iu_gpr_10__5_), .Y(_6564_) );
	OAI21X1 OAI21X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf1), .B(_6558__bF_buf4), .C(_6564_), .Y(_2273_) );
	OAI21X1 OAI21X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2590__bF_buf0), .C(csr_gpr_iu_gpr_10__6_), .Y(_6565_) );
	OAI21X1 OAI21X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf1), .B(_6558__bF_buf3), .C(_6565_), .Y(_2274_) );
	OAI21X1 OAI21X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2590__bF_buf12), .C(csr_gpr_iu_gpr_10__7_), .Y(_6566_) );
	OAI21X1 OAI21X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf1), .B(_6558__bF_buf2), .C(_6566_), .Y(_2275_) );
	OAI21X1 OAI21X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2590__bF_buf11), .C(csr_gpr_iu_gpr_10__8_), .Y(_6567_) );
	OAI21X1 OAI21X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf1), .B(_6558__bF_buf1), .C(_6567_), .Y(_2276_) );
	OAI21X1 OAI21X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2590__bF_buf10), .C(csr_gpr_iu_gpr_10__9_), .Y(_6568_) );
	OAI21X1 OAI21X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf1), .B(_6558__bF_buf0), .C(_6568_), .Y(_2277_) );
	OAI21X1 OAI21X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2590__bF_buf9), .C(csr_gpr_iu_gpr_10__10_), .Y(_6569_) );
	OAI21X1 OAI21X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf1), .B(_6558__bF_buf4), .C(_6569_), .Y(_2278_) );
	OAI21X1 OAI21X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2590__bF_buf8), .C(csr_gpr_iu_gpr_10__11_), .Y(_6570_) );
	OAI21X1 OAI21X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf1), .B(_6558__bF_buf3), .C(_6570_), .Y(_2279_) );
	OAI21X1 OAI21X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2590__bF_buf7), .C(csr_gpr_iu_gpr_10__12_), .Y(_6571_) );
	OAI21X1 OAI21X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf1), .B(_6558__bF_buf2), .C(_6571_), .Y(_2280_) );
	OAI21X1 OAI21X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_10__13_), .Y(_6572_) );
	OAI21X1 OAI21X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf1), .B(_6558__bF_buf1), .C(_6572_), .Y(_2281_) );
	OAI21X1 OAI21X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2590__bF_buf5), .C(csr_gpr_iu_gpr_10__14_), .Y(_6573_) );
	OAI21X1 OAI21X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf1), .B(_6558__bF_buf0), .C(_6573_), .Y(_2282_) );
	OAI21X1 OAI21X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2590__bF_buf4), .C(csr_gpr_iu_gpr_10__15_), .Y(_6574_) );
	OAI21X1 OAI21X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf1), .B(_6558__bF_buf4), .C(_6574_), .Y(_2283_) );
	OAI21X1 OAI21X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2590__bF_buf3), .C(csr_gpr_iu_gpr_10__16_), .Y(_6575_) );
	OAI21X1 OAI21X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf1), .B(_6558__bF_buf3), .C(_6575_), .Y(_2284_) );
	OAI21X1 OAI21X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2590__bF_buf2), .C(csr_gpr_iu_gpr_10__17_), .Y(_6576_) );
	OAI21X1 OAI21X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf1), .B(_6558__bF_buf2), .C(_6576_), .Y(_2285_) );
	OAI21X1 OAI21X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2590__bF_buf1), .C(csr_gpr_iu_gpr_10__18_), .Y(_6577_) );
	OAI21X1 OAI21X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf1), .B(_6558__bF_buf1), .C(_6577_), .Y(_2286_) );
	OAI21X1 OAI21X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2590__bF_buf0), .C(csr_gpr_iu_gpr_10__19_), .Y(_6578_) );
	OAI21X1 OAI21X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf1), .B(_6558__bF_buf0), .C(_6578_), .Y(_2287_) );
	OAI21X1 OAI21X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2590__bF_buf12), .C(csr_gpr_iu_gpr_10__20_), .Y(_6579_) );
	OAI21X1 OAI21X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf1), .B(_6558__bF_buf4), .C(_6579_), .Y(_2288_) );
	OAI21X1 OAI21X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2590__bF_buf11), .C(csr_gpr_iu_gpr_10__21_), .Y(_6580_) );
	OAI21X1 OAI21X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf1), .B(_6558__bF_buf3), .C(_6580_), .Y(_2289_) );
	OAI21X1 OAI21X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf1), .B(_2590__bF_buf10), .C(csr_gpr_iu_gpr_10__22_), .Y(_6581_) );
	OAI21X1 OAI21X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf1), .B(_6558__bF_buf2), .C(_6581_), .Y(_2290_) );
	OAI21X1 OAI21X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf0), .B(_2590__bF_buf9), .C(csr_gpr_iu_gpr_10__23_), .Y(_6582_) );
	OAI21X1 OAI21X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf1), .B(_6558__bF_buf1), .C(_6582_), .Y(_2291_) );
	OAI21X1 OAI21X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf10), .B(_2590__bF_buf8), .C(csr_gpr_iu_gpr_10__24_), .Y(_6583_) );
	OAI21X1 OAI21X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf1), .B(_6558__bF_buf0), .C(_6583_), .Y(_2292_) );
	OAI21X1 OAI21X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf9), .B(_2590__bF_buf7), .C(csr_gpr_iu_gpr_10__25_), .Y(_6584_) );
	OAI21X1 OAI21X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf1), .B(_6558__bF_buf4), .C(_6584_), .Y(_2293_) );
	OAI21X1 OAI21X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf8), .B(_2590__bF_buf6), .C(csr_gpr_iu_gpr_10__26_), .Y(_6585_) );
	OAI21X1 OAI21X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf1), .B(_6558__bF_buf3), .C(_6585_), .Y(_2294_) );
	OAI21X1 OAI21X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf7), .B(_2590__bF_buf5), .C(csr_gpr_iu_gpr_10__27_), .Y(_6586_) );
	OAI21X1 OAI21X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf1), .B(_6558__bF_buf2), .C(_6586_), .Y(_2295_) );
	OAI21X1 OAI21X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf6), .B(_2590__bF_buf4), .C(csr_gpr_iu_gpr_10__28_), .Y(_6587_) );
	OAI21X1 OAI21X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf1), .B(_6558__bF_buf1), .C(_6587_), .Y(_2296_) );
	OAI21X1 OAI21X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf5), .B(_2590__bF_buf3), .C(csr_gpr_iu_gpr_10__29_), .Y(_6588_) );
	OAI21X1 OAI21X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf1), .B(_6558__bF_buf0), .C(_6588_), .Y(_2297_) );
	OAI21X1 OAI21X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf4), .B(_2590__bF_buf2), .C(csr_gpr_iu_gpr_10__30_), .Y(_6589_) );
	OAI21X1 OAI21X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_6558__bF_buf4), .C(_6589_), .Y(_2298_) );
	OAI21X1 OAI21X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf3), .B(_2590__bF_buf1), .C(csr_gpr_iu_gpr_10__31_), .Y(_6590_) );
	OAI21X1 OAI21X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf1), .B(_6558__bF_buf3), .C(_6590_), .Y(_2299_) );
	OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_6426__bF_buf2), .B(_2625__bF_buf1), .Y(_6591_) );
	OAI21X1 OAI21X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6426__bF_buf1), .C(csr_gpr_iu_gpr_11__0_), .Y(_6592_) );
	OAI21X1 OAI21X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_2460__bF_buf0), .B(_6591__bF_buf4), .C(_6592_), .Y(_2300_) );
	OAI21X1 OAI21X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6426__bF_buf0), .C(csr_gpr_iu_gpr_11__1_), .Y(_6593_) );
	OAI21X1 OAI21X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_2489__bF_buf0), .B(_6591__bF_buf3), .C(_6593_), .Y(_2301_) );
	OAI21X1 OAI21X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6426__bF_buf10), .C(csr_gpr_iu_gpr_11__2_), .Y(_6594_) );
	OAI21X1 OAI21X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_2491__bF_buf0), .B(_6591__bF_buf2), .C(_6594_), .Y(_2302_) );
	OAI21X1 OAI21X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6426__bF_buf9), .C(csr_gpr_iu_gpr_11__3_), .Y(_6595_) );
	OAI21X1 OAI21X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_2493__bF_buf0), .B(_6591__bF_buf1), .C(_6595_), .Y(_2303_) );
	OAI21X1 OAI21X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6426__bF_buf8), .C(csr_gpr_iu_gpr_11__4_), .Y(_6596_) );
	OAI21X1 OAI21X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_2495__bF_buf0), .B(_6591__bF_buf0), .C(_6596_), .Y(_2304_) );
	OAI21X1 OAI21X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6426__bF_buf7), .C(csr_gpr_iu_gpr_11__5_), .Y(_6597_) );
	OAI21X1 OAI21X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_2497__bF_buf0), .B(_6591__bF_buf4), .C(_6597_), .Y(_2305_) );
	OAI21X1 OAI21X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6426__bF_buf6), .C(csr_gpr_iu_gpr_11__6_), .Y(_6598_) );
	OAI21X1 OAI21X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_2499__bF_buf0), .B(_6591__bF_buf3), .C(_6598_), .Y(_2306_) );
	OAI21X1 OAI21X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6426__bF_buf5), .C(csr_gpr_iu_gpr_11__7_), .Y(_6599_) );
	OAI21X1 OAI21X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_2501__bF_buf0), .B(_6591__bF_buf2), .C(_6599_), .Y(_2307_) );
	OAI21X1 OAI21X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6426__bF_buf4), .C(csr_gpr_iu_gpr_11__8_), .Y(_6600_) );
	OAI21X1 OAI21X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_2503__bF_buf0), .B(_6591__bF_buf1), .C(_6600_), .Y(_2308_) );
	OAI21X1 OAI21X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6426__bF_buf3), .C(csr_gpr_iu_gpr_11__9_), .Y(_6601_) );
	OAI21X1 OAI21X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_2505__bF_buf0), .B(_6591__bF_buf0), .C(_6601_), .Y(_2309_) );
	OAI21X1 OAI21X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6426__bF_buf2), .C(csr_gpr_iu_gpr_11__10_), .Y(_6602_) );
	OAI21X1 OAI21X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_2507__bF_buf0), .B(_6591__bF_buf4), .C(_6602_), .Y(_2310_) );
	OAI21X1 OAI21X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6426__bF_buf1), .C(csr_gpr_iu_gpr_11__11_), .Y(_6603_) );
	OAI21X1 OAI21X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_2509__bF_buf0), .B(_6591__bF_buf3), .C(_6603_), .Y(_2311_) );
	OAI21X1 OAI21X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6426__bF_buf0), .C(csr_gpr_iu_gpr_11__12_), .Y(_6604_) );
	OAI21X1 OAI21X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_2511__bF_buf0), .B(_6591__bF_buf2), .C(_6604_), .Y(_2312_) );
	OAI21X1 OAI21X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6426__bF_buf10), .C(csr_gpr_iu_gpr_11__13_), .Y(_6605_) );
	OAI21X1 OAI21X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_2513__bF_buf0), .B(_6591__bF_buf1), .C(_6605_), .Y(_2313_) );
	OAI21X1 OAI21X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6426__bF_buf9), .C(csr_gpr_iu_gpr_11__14_), .Y(_6606_) );
	OAI21X1 OAI21X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_2515__bF_buf0), .B(_6591__bF_buf0), .C(_6606_), .Y(_2314_) );
	OAI21X1 OAI21X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6426__bF_buf8), .C(csr_gpr_iu_gpr_11__15_), .Y(_6607_) );
	OAI21X1 OAI21X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_2517__bF_buf0), .B(_6591__bF_buf4), .C(_6607_), .Y(_2315_) );
	OAI21X1 OAI21X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6426__bF_buf7), .C(csr_gpr_iu_gpr_11__16_), .Y(_6608_) );
	OAI21X1 OAI21X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_2519__bF_buf0), .B(_6591__bF_buf3), .C(_6608_), .Y(_2316_) );
	OAI21X1 OAI21X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf13), .B(_6426__bF_buf6), .C(csr_gpr_iu_gpr_11__17_), .Y(_6609_) );
	OAI21X1 OAI21X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_2521__bF_buf0), .B(_6591__bF_buf2), .C(_6609_), .Y(_2317_) );
	OAI21X1 OAI21X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf12), .B(_6426__bF_buf5), .C(csr_gpr_iu_gpr_11__18_), .Y(_6610_) );
	OAI21X1 OAI21X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_2523__bF_buf0), .B(_6591__bF_buf1), .C(_6610_), .Y(_2318_) );
	OAI21X1 OAI21X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf11), .B(_6426__bF_buf4), .C(csr_gpr_iu_gpr_11__19_), .Y(_6611_) );
	OAI21X1 OAI21X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_2525__bF_buf0), .B(_6591__bF_buf0), .C(_6611_), .Y(_2319_) );
	OAI21X1 OAI21X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf10), .B(_6426__bF_buf3), .C(csr_gpr_iu_gpr_11__20_), .Y(_6612_) );
	OAI21X1 OAI21X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_2527__bF_buf0), .B(_6591__bF_buf4), .C(_6612_), .Y(_2320_) );
	OAI21X1 OAI21X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf9), .B(_6426__bF_buf2), .C(csr_gpr_iu_gpr_11__21_), .Y(_6613_) );
	OAI21X1 OAI21X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_2529__bF_buf0), .B(_6591__bF_buf3), .C(_6613_), .Y(_2321_) );
	OAI21X1 OAI21X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf8), .B(_6426__bF_buf1), .C(csr_gpr_iu_gpr_11__22_), .Y(_6614_) );
	OAI21X1 OAI21X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_2531__bF_buf0), .B(_6591__bF_buf2), .C(_6614_), .Y(_2322_) );
	OAI21X1 OAI21X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf7), .B(_6426__bF_buf0), .C(csr_gpr_iu_gpr_11__23_), .Y(_6615_) );
	OAI21X1 OAI21X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_2533__bF_buf0), .B(_6591__bF_buf1), .C(_6615_), .Y(_2323_) );
	OAI21X1 OAI21X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf6), .B(_6426__bF_buf10), .C(csr_gpr_iu_gpr_11__24_), .Y(_6616_) );
	OAI21X1 OAI21X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_2535__bF_buf0), .B(_6591__bF_buf0), .C(_6616_), .Y(_2324_) );
	OAI21X1 OAI21X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf5), .B(_6426__bF_buf9), .C(csr_gpr_iu_gpr_11__25_), .Y(_6617_) );
	OAI21X1 OAI21X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_2537__bF_buf0), .B(_6591__bF_buf4), .C(_6617_), .Y(_2325_) );
	OAI21X1 OAI21X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf4), .B(_6426__bF_buf8), .C(csr_gpr_iu_gpr_11__26_), .Y(_6618_) );
	OAI21X1 OAI21X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_2539__bF_buf0), .B(_6591__bF_buf3), .C(_6618_), .Y(_2326_) );
	OAI21X1 OAI21X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf3), .B(_6426__bF_buf7), .C(csr_gpr_iu_gpr_11__27_), .Y(_6619_) );
	OAI21X1 OAI21X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_2541__bF_buf0), .B(_6591__bF_buf2), .C(_6619_), .Y(_2327_) );
	OAI21X1 OAI21X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf2), .B(_6426__bF_buf6), .C(csr_gpr_iu_gpr_11__28_), .Y(_6620_) );
	OAI21X1 OAI21X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_2543__bF_buf0), .B(_6591__bF_buf1), .C(_6620_), .Y(_2328_) );
	OAI21X1 OAI21X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf1), .B(_6426__bF_buf5), .C(csr_gpr_iu_gpr_11__29_), .Y(_6621_) );
	OAI21X1 OAI21X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_2545__bF_buf0), .B(_6591__bF_buf0), .C(_6621_), .Y(_2329_) );
	OAI21X1 OAI21X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf0), .B(_6426__bF_buf4), .C(csr_gpr_iu_gpr_11__30_), .Y(_6622_) );
	OAI21X1 OAI21X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_6591__bF_buf4), .C(_6622_), .Y(_2330_) );
	OAI21X1 OAI21X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_2625__bF_buf14), .B(_6426__bF_buf3), .C(csr_gpr_iu_gpr_11__31_), .Y(_6623_) );
	OAI21X1 OAI21X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_2549__bF_buf0), .B(_6591__bF_buf3), .C(_6623_), .Y(_2331_) );
	NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_st_page_fault_reg), .B(biu_exce_chk_st_page_fault), .Y(_6624_) );
	INVX1 INVX1_1113 ( .gnd(gnd), .vdd(vdd), .A(_6624_), .Y(csr_gpr_iu_int_ctrl_st_page_fault) );
	NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_reg), .B(biu_exce_chk_ins_page_fault), .Y(_6625_) );
	INVX8 INVX8_53 ( .gnd(gnd), .vdd(vdd), .A(_6625_), .Y(csr_gpr_iu_ins_page_fault) );
	NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ld_page_fault_reg), .B(biu_exce_chk_ld_page_fault), .Y(_6626_) );
	INVX1 INVX1_1114 ( .gnd(gnd), .vdd(vdd), .A(_6626_), .Y(csr_gpr_iu_int_ctrl_ld_page_fault) );
	OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_addr_mis_reg), .B(biu_exce_chk_ins_addr_mis), .Y(csr_gpr_iu_ins_addr_mis) );
	OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_acc_fault_reg), .B(biu_exce_chk_ins_acc_fault), .Y(csr_gpr_iu_ins_acc_fault) );
	NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_load_addr_mis_reg), .B(biu_exce_chk_load_addr_mis), .Y(_6627_) );
	INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .Y(csr_gpr_iu_int_ctrl_load_addr_mis) );
	NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_load_acc_fault_reg), .B(biu_exce_chk_load_acc_fault), .Y(_6628_) );
	INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_6628_), .Y(csr_gpr_iu_int_ctrl_load_acc_fault) );
	NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_st_addr_mis_reg), .B(biu_exce_chk_st_addr_mis), .Y(_6629_) );
	INVX1 INVX1_1115 ( .gnd(gnd), .vdd(vdd), .A(_6629_), .Y(csr_gpr_iu_int_ctrl_st_addr_mis) );
	NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_st_acc_fault_reg), .B(biu_exce_chk_st_acc_fault), .Y(_6630_) );
	INVX1 INVX1_1116 ( .gnd(gnd), .vdd(vdd), .A(_6630_), .Y(csr_gpr_iu_int_ctrl_st_acc_fault) );
	NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_6628_), .B(_6629_), .C(_6630_), .Y(_6631_) );
	INVX1 INVX1_1117 ( .gnd(gnd), .vdd(vdd), .A(_6631_), .Y(_6632_) );
	NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_addr_mis), .B(csr_gpr_iu_ins_acc_fault), .Y(_6633_) );
	NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_6624_), .B(_6625_), .Y(_6634_) );
	NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_6626_), .B(_6627_), .Y(_6635_) );
	NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_6634_), .B(_6635_), .Y(_6636_) );
	NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_6633_), .B(_6632_), .C(_6636_), .Y(_6637_) );
	OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(biu_rdy_biu), .Y(_6638_) );
	INVX1 INVX1_1118 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .Y(_6639_) );
	INVX1 INVX1_1119 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .Y(_6640_) );
	INVX1 INVX1_1120 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .Y(_6641_) );
	NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_6640_), .B(_6641_), .Y(_6642_) );
	NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_6642_), .B(_6639_), .Y(_6643_) );
	NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(_6641_), .Y(_6644_) );
	NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(_6644_), .Y(_6645_) );
	OAI22X1 OAI22X1_643 ( .gnd(gnd), .vdd(vdd), .A(_6643_), .B(_6645_), .C(_6638_), .D(_6637_), .Y(_6646_) );
	NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_6640_), .B(biu_exce_chk_statu_cpu_0_), .C(_2465_), .Y(_6647_) );
	INVX1 INVX1_1121 ( .gnd(gnd), .vdd(vdd), .A(_6647_), .Y(_6648_) );
	NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ebreak), .B(csr_gpr_iu_ecall), .C(csr_gpr_iu_ill_ins), .Y(_6649_) );
	NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_ins_flow_3_), .B(csr_gpr_iu_ins_dec_ins_flow_3_), .Y(_6650_) );
	AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rdy_exu), .B(csr_gpr_iu_ins_dec_ins_flow_1_), .Y(_6651_) );
	NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_6650_), .B(_6651_), .Y(_6652_) );
	NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_6641_), .B(_6652_), .Y(_6653_) );
	AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rdy_exu), .B(csr_gpr_iu_ins_dec_ins_flow_0_), .Y(_6654_) );
	NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_6650_), .B(_6654_), .Y(_6655_) );
	NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_6655_), .B(_6653_), .Y(_6656_) );
	NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_6656_), .Y(_6657_) );
	INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_acc), .Y(_6658_) );
	NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(_2467_), .Y(_6659_) );
	NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_2_), .C(_2467_), .Y(_6660_) );
	NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(_6659_), .C(_6660_), .Y(_6661_) );
	OAI21X1 OAI21X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_6659_), .C(_6661_), .Y(_6662_) );
	NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(_6640_), .Y(_6663_) );
	INVX1 INVX1_1122 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .Y(_6664_) );
	NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(_6664_), .Y(_6665_) );
	NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_6663_), .B(_6665_), .Y(_6666_) );
	AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(csr_gpr_iu_rdy_exu), .C(_6648_), .Y(_6667_) );
	AOI22X1 AOI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_6662_), .B(_6667_), .C(_6648_), .D(_6657_), .Y(_6668_) );
	AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_6668_), .B(_6646_), .C(rst_bF_buf69), .Y(_1467__0_) );
	NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(_6659_), .C(_6660_), .Y(_6669_) );
	OAI21X1 OAI21X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_6659_), .C(_6669_), .Y(_6670_) );
	NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rdy_exu), .B(_6666_), .Y(_6671_) );
	OAI21X1 OAI21X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6665_), .C(_6671_), .Y(_6672_) );
	NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6665_), .Y(_6673_) );
	OAI21X1 OAI21X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_6640_), .B(biu_rdy_biu), .C(_6673_), .Y(_6674_) );
	OAI22X1 OAI22X1_644 ( .gnd(gnd), .vdd(vdd), .A(_6637_), .B(_6674_), .C(_6672_), .D(_6670_), .Y(_6675_) );
	NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_6643_), .B(_6637_), .Y(_6676_) );
	INVX1 INVX1_1123 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_ins_flow_0_), .Y(_6677_) );
	NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6652_), .Y(_6678_) );
	INVX1 INVX1_1124 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_ins_flow_1_), .Y(_6679_) );
	NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_6679_), .B(_6650_), .C(_6654_), .Y(_6680_) );
	NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6650_), .C(_6651_), .Y(_6681_) );
	NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_6680_), .C(_6681_), .Y(_6682_) );
	OAI21X1 OAI21X1_3160 ( .gnd(gnd), .vdd(vdd), .A(_6678_), .B(_6682_), .C(_6648_), .Y(_6683_) );
	AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_6676_), .B(_6683_), .Y(_6684_) );
	AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_6684_), .B(_6675_), .C(rst_bF_buf68), .Y(_1467__1_) );
	NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_6659_), .Y(_6685_) );
	NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_6647_), .Y(_6686_) );
	NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_6686_), .B(_6685_), .Y(_6687_) );
	AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_6676_), .B(_6687_), .Y(_6688_) );
	NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(_2467_), .Y(_6689_) );
	AOI22X1 AOI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(_6689_), .C(_6645_), .D(_6637_), .Y(_6690_) );
	AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_6688_), .B(_6690_), .C(rst_bF_buf67), .Y(_1467__2_) );
	INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf66), .Y(_6691_) );
	NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6639_), .Y(_6692_) );
	NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(biu_rdy_biu), .B(_6664_), .Y(_6693_) );
	OAI21X1 OAI21X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .B(_6637_), .C(_6692_), .Y(_6694_) );
	NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rdy_exu), .B(csr_gpr_iu_ins_dec_ins_flow_0_), .C(csr_gpr_iu_ins_dec_ins_flow_1_), .Y(_6695_) );
	INVX1 INVX1_1125 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .Y(_6696_) );
	AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_6696_), .B(_6650_), .C(biu_exce_chk_statu_cpu_3_), .Y(_6697_) );
	OAI21X1 OAI21X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_6697_), .B(_6682_), .C(_6649_), .Y(_6698_) );
	NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_6648_), .B(_6698_), .Y(_6699_) );
	OAI21X1 OAI21X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_6664_), .B(_2466_), .C(biu_exce_chk_statu_cpu_3_), .Y(_6700_) );
	OAI21X1 OAI21X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_6659_), .C(_6700_), .Y(_6701_) );
	AOI22X1 AOI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_6671_), .B(_6701_), .C(_6643_), .D(_6637_), .Y(_6702_) );
	NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_6702_), .B(_6694_), .C(_6699_), .Y(_6703_) );
	AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_6703_), .B(_6691_), .Y(_1467__3_) );
	AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_st_page_fault), .Y(_1466_) );
	AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_ld_page_fault), .Y(_1461_) );
	AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_ins_page_fault), .Y(_1460_) );
	AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_st_acc_fault), .Y(_1464_) );
	AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_st_addr_mis), .Y(_1465_) );
	AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_load_acc_fault), .Y(_1462_) );
	AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_load_addr_mis), .Y(_1463_) );
	AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_ins_acc_fault), .Y(_1458_) );
	AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(biu_exce_chk_ins_addr_mis), .Y(_1459_) );
	DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_2332_), .Q(csr_gpr_iu_gpr_29__0_) );
	DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_2333_), .Q(csr_gpr_iu_gpr_29__1_) );
	DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_2334_), .Q(csr_gpr_iu_gpr_29__2_) );
	DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_2335_), .Q(csr_gpr_iu_gpr_29__3_) );
	DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_2336_), .Q(csr_gpr_iu_gpr_29__4_) );
	DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_2337_), .Q(csr_gpr_iu_gpr_29__5_) );
	DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_2338_), .Q(csr_gpr_iu_gpr_29__6_) );
	DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_2339_), .Q(csr_gpr_iu_gpr_29__7_) );
	DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_2340_), .Q(csr_gpr_iu_gpr_29__8_) );
	DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_2341_), .Q(csr_gpr_iu_gpr_29__9_) );
	DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_2342_), .Q(csr_gpr_iu_gpr_29__10_) );
	DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_2343_), .Q(csr_gpr_iu_gpr_29__11_) );
	DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_2344_), .Q(csr_gpr_iu_gpr_29__12_) );
	DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_2345_), .Q(csr_gpr_iu_gpr_29__13_) );
	DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_2346_), .Q(csr_gpr_iu_gpr_29__14_) );
	DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_2347_), .Q(csr_gpr_iu_gpr_29__15_) );
	DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_2348_), .Q(csr_gpr_iu_gpr_29__16_) );
	DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_2349_), .Q(csr_gpr_iu_gpr_29__17_) );
	DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_2350_), .Q(csr_gpr_iu_gpr_29__18_) );
	DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_2351_), .Q(csr_gpr_iu_gpr_29__19_) );
	DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_2352_), .Q(csr_gpr_iu_gpr_29__20_) );
	DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_2353_), .Q(csr_gpr_iu_gpr_29__21_) );
	DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_2354_), .Q(csr_gpr_iu_gpr_29__22_) );
	DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_2355_), .Q(csr_gpr_iu_gpr_29__23_) );
	DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_2356_), .Q(csr_gpr_iu_gpr_29__24_) );
	DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_2357_), .Q(csr_gpr_iu_gpr_29__25_) );
	DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_2358_), .Q(csr_gpr_iu_gpr_29__26_) );
	DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_2359_), .Q(csr_gpr_iu_gpr_29__27_) );
	DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_2360_), .Q(csr_gpr_iu_gpr_29__28_) );
	DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_2361_), .Q(csr_gpr_iu_gpr_29__29_) );
	DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_2362_), .Q(csr_gpr_iu_gpr_29__30_) );
	DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_2363_), .Q(csr_gpr_iu_gpr_29__31_) );
	DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_2428_), .Q(csr_gpr_iu_gpr_27__0_) );
	DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_2429_), .Q(csr_gpr_iu_gpr_27__1_) );
	DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_2430_), .Q(csr_gpr_iu_gpr_27__2_) );
	DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_2431_), .Q(csr_gpr_iu_gpr_27__3_) );
	DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_2432_), .Q(csr_gpr_iu_gpr_27__4_) );
	DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_2433_), .Q(csr_gpr_iu_gpr_27__5_) );
	DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_2434_), .Q(csr_gpr_iu_gpr_27__6_) );
	DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_2435_), .Q(csr_gpr_iu_gpr_27__7_) );
	DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_2436_), .Q(csr_gpr_iu_gpr_27__8_) );
	DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_2437_), .Q(csr_gpr_iu_gpr_27__9_) );
	DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_2438_), .Q(csr_gpr_iu_gpr_27__10_) );
	DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_2439_), .Q(csr_gpr_iu_gpr_27__11_) );
	DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_2440_), .Q(csr_gpr_iu_gpr_27__12_) );
	DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_2441_), .Q(csr_gpr_iu_gpr_27__13_) );
	DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_2442_), .Q(csr_gpr_iu_gpr_27__14_) );
	DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_2443_), .Q(csr_gpr_iu_gpr_27__15_) );
	DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_2444_), .Q(csr_gpr_iu_gpr_27__16_) );
	DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_2445_), .Q(csr_gpr_iu_gpr_27__17_) );
	DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_2446_), .Q(csr_gpr_iu_gpr_27__18_) );
	DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_2447_), .Q(csr_gpr_iu_gpr_27__19_) );
	DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_2448_), .Q(csr_gpr_iu_gpr_27__20_) );
	DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_2449_), .Q(csr_gpr_iu_gpr_27__21_) );
	DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_2450_), .Q(csr_gpr_iu_gpr_27__22_) );
	DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_2451_), .Q(csr_gpr_iu_gpr_27__23_) );
	DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_2452_), .Q(csr_gpr_iu_gpr_27__24_) );
	DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_2453_), .Q(csr_gpr_iu_gpr_27__25_) );
	DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_2454_), .Q(csr_gpr_iu_gpr_27__26_) );
	DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_2455_), .Q(csr_gpr_iu_gpr_27__27_) );
	DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_2456_), .Q(csr_gpr_iu_gpr_27__28_) );
	DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_2457_), .Q(csr_gpr_iu_gpr_27__29_) );
	DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_2458_), .Q(csr_gpr_iu_gpr_27__30_) );
	DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_2459_), .Q(csr_gpr_iu_gpr_27__31_) );
	DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1628_), .Q(csr_gpr_iu_gpr_23__0_) );
	DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1629_), .Q(csr_gpr_iu_gpr_23__1_) );
	DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1630_), .Q(csr_gpr_iu_gpr_23__2_) );
	DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1631_), .Q(csr_gpr_iu_gpr_23__3_) );
	DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1632_), .Q(csr_gpr_iu_gpr_23__4_) );
	DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1633_), .Q(csr_gpr_iu_gpr_23__5_) );
	DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1634_), .Q(csr_gpr_iu_gpr_23__6_) );
	DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1635_), .Q(csr_gpr_iu_gpr_23__7_) );
	DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1636_), .Q(csr_gpr_iu_gpr_23__8_) );
	DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1637_), .Q(csr_gpr_iu_gpr_23__9_) );
	DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1638_), .Q(csr_gpr_iu_gpr_23__10_) );
	DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1639_), .Q(csr_gpr_iu_gpr_23__11_) );
	DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1640_), .Q(csr_gpr_iu_gpr_23__12_) );
	DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1641_), .Q(csr_gpr_iu_gpr_23__13_) );
	DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1642_), .Q(csr_gpr_iu_gpr_23__14_) );
	DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1643_), .Q(csr_gpr_iu_gpr_23__15_) );
	DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1644_), .Q(csr_gpr_iu_gpr_23__16_) );
	DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1645_), .Q(csr_gpr_iu_gpr_23__17_) );
	DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1646_), .Q(csr_gpr_iu_gpr_23__18_) );
	DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1647_), .Q(csr_gpr_iu_gpr_23__19_) );
	DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1648_), .Q(csr_gpr_iu_gpr_23__20_) );
	DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1649_), .Q(csr_gpr_iu_gpr_23__21_) );
	DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1650_), .Q(csr_gpr_iu_gpr_23__22_) );
	DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1651_), .Q(csr_gpr_iu_gpr_23__23_) );
	DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1652_), .Q(csr_gpr_iu_gpr_23__24_) );
	DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1653_), .Q(csr_gpr_iu_gpr_23__25_) );
	DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1654_), .Q(csr_gpr_iu_gpr_23__26_) );
	DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1655_), .Q(csr_gpr_iu_gpr_23__27_) );
	DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1656_), .Q(csr_gpr_iu_gpr_23__28_) );
	DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1657_), .Q(csr_gpr_iu_gpr_23__29_) );
	DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_1658_), .Q(csr_gpr_iu_gpr_23__30_) );
	DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_1659_), .Q(csr_gpr_iu_gpr_23__31_) );
	DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_1692_), .Q(csr_gpr_iu_gpr_18__0_) );
	DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1693_), .Q(csr_gpr_iu_gpr_18__1_) );
	DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_1694_), .Q(csr_gpr_iu_gpr_18__2_) );
	DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_1695_), .Q(csr_gpr_iu_gpr_18__3_) );
	DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_1696_), .Q(csr_gpr_iu_gpr_18__4_) );
	DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_1697_), .Q(csr_gpr_iu_gpr_18__5_) );
	DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_1698_), .Q(csr_gpr_iu_gpr_18__6_) );
	DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_1699_), .Q(csr_gpr_iu_gpr_18__7_) );
	DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_1700_), .Q(csr_gpr_iu_gpr_18__8_) );
	DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_1701_), .Q(csr_gpr_iu_gpr_18__9_) );
	DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_1702_), .Q(csr_gpr_iu_gpr_18__10_) );
	DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_1703_), .Q(csr_gpr_iu_gpr_18__11_) );
	DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_1704_), .Q(csr_gpr_iu_gpr_18__12_) );
	DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_1705_), .Q(csr_gpr_iu_gpr_18__13_) );
	DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_1706_), .Q(csr_gpr_iu_gpr_18__14_) );
	DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_1707_), .Q(csr_gpr_iu_gpr_18__15_) );
	DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_1708_), .Q(csr_gpr_iu_gpr_18__16_) );
	DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_1709_), .Q(csr_gpr_iu_gpr_18__17_) );
	DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_1710_), .Q(csr_gpr_iu_gpr_18__18_) );
	DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_1711_), .Q(csr_gpr_iu_gpr_18__19_) );
	DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_1712_), .Q(csr_gpr_iu_gpr_18__20_) );
	DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_1713_), .Q(csr_gpr_iu_gpr_18__21_) );
	DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_1714_), .Q(csr_gpr_iu_gpr_18__22_) );
	DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_1715_), .Q(csr_gpr_iu_gpr_18__23_) );
	DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_1716_), .Q(csr_gpr_iu_gpr_18__24_) );
	DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_1717_), .Q(csr_gpr_iu_gpr_18__25_) );
	DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1718_), .Q(csr_gpr_iu_gpr_18__26_) );
	DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_1719_), .Q(csr_gpr_iu_gpr_18__27_) );
	DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_1720_), .Q(csr_gpr_iu_gpr_18__28_) );
	DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_1721_), .Q(csr_gpr_iu_gpr_18__29_) );
	DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_1722_), .Q(csr_gpr_iu_gpr_18__30_) );
	DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_1723_), .Q(csr_gpr_iu_gpr_18__31_) );
	DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_2396_), .Q(csr_gpr_iu_gpr_26__0_) );
	DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_2397_), .Q(csr_gpr_iu_gpr_26__1_) );
	DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_2398_), .Q(csr_gpr_iu_gpr_26__2_) );
	DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_2399_), .Q(csr_gpr_iu_gpr_26__3_) );
	DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_2400_), .Q(csr_gpr_iu_gpr_26__4_) );
	DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_2401_), .Q(csr_gpr_iu_gpr_26__5_) );
	DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_2402_), .Q(csr_gpr_iu_gpr_26__6_) );
	DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_2403_), .Q(csr_gpr_iu_gpr_26__7_) );
	DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_2404_), .Q(csr_gpr_iu_gpr_26__8_) );
	DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2405_), .Q(csr_gpr_iu_gpr_26__9_) );
	DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_2406_), .Q(csr_gpr_iu_gpr_26__10_) );
	DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_2407_), .Q(csr_gpr_iu_gpr_26__11_) );
	DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_2408_), .Q(csr_gpr_iu_gpr_26__12_) );
	DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_2409_), .Q(csr_gpr_iu_gpr_26__13_) );
	DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2410_), .Q(csr_gpr_iu_gpr_26__14_) );
	DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2411_), .Q(csr_gpr_iu_gpr_26__15_) );
	DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2412_), .Q(csr_gpr_iu_gpr_26__16_) );
	DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2413_), .Q(csr_gpr_iu_gpr_26__17_) );
	DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2414_), .Q(csr_gpr_iu_gpr_26__18_) );
	DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2415_), .Q(csr_gpr_iu_gpr_26__19_) );
	DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2416_), .Q(csr_gpr_iu_gpr_26__20_) );
	DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2417_), .Q(csr_gpr_iu_gpr_26__21_) );
	DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_2418_), .Q(csr_gpr_iu_gpr_26__22_) );
	DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_2419_), .Q(csr_gpr_iu_gpr_26__23_) );
	DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_2420_), .Q(csr_gpr_iu_gpr_26__24_) );
	DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_2421_), .Q(csr_gpr_iu_gpr_26__25_) );
	DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_2422_), .Q(csr_gpr_iu_gpr_26__26_) );
	DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_2423_), .Q(csr_gpr_iu_gpr_26__27_) );
	DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_2424_), .Q(csr_gpr_iu_gpr_26__28_) );
	DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_2425_), .Q(csr_gpr_iu_gpr_26__29_) );
	DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_2426_), .Q(csr_gpr_iu_gpr_26__30_) );
	DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_2427_), .Q(csr_gpr_iu_gpr_26__31_) );
	DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_1564_), .Q(csr_gpr_iu_gpr_21__0_) );
	DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_1565_), .Q(csr_gpr_iu_gpr_21__1_) );
	DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_1566_), .Q(csr_gpr_iu_gpr_21__2_) );
	DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_1567_), .Q(csr_gpr_iu_gpr_21__3_) );
	DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_1568_), .Q(csr_gpr_iu_gpr_21__4_) );
	DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_1569_), .Q(csr_gpr_iu_gpr_21__5_) );
	DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_1570_), .Q(csr_gpr_iu_gpr_21__6_) );
	DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_1571_), .Q(csr_gpr_iu_gpr_21__7_) );
	DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_1572_), .Q(csr_gpr_iu_gpr_21__8_) );
	DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_1573_), .Q(csr_gpr_iu_gpr_21__9_) );
	DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_1574_), .Q(csr_gpr_iu_gpr_21__10_) );
	DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_1575_), .Q(csr_gpr_iu_gpr_21__11_) );
	DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_1576_), .Q(csr_gpr_iu_gpr_21__12_) );
	DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_1577_), .Q(csr_gpr_iu_gpr_21__13_) );
	DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_1578_), .Q(csr_gpr_iu_gpr_21__14_) );
	DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_1579_), .Q(csr_gpr_iu_gpr_21__15_) );
	DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_1580_), .Q(csr_gpr_iu_gpr_21__16_) );
	DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_1581_), .Q(csr_gpr_iu_gpr_21__17_) );
	DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_1582_), .Q(csr_gpr_iu_gpr_21__18_) );
	DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_1583_), .Q(csr_gpr_iu_gpr_21__19_) );
	DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_1584_), .Q(csr_gpr_iu_gpr_21__20_) );
	DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_1585_), .Q(csr_gpr_iu_gpr_21__21_) );
	DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_1586_), .Q(csr_gpr_iu_gpr_21__22_) );
	DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_1587_), .Q(csr_gpr_iu_gpr_21__23_) );
	DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_1588_), .Q(csr_gpr_iu_gpr_21__24_) );
	DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_1589_), .Q(csr_gpr_iu_gpr_21__25_) );
	DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_1590_), .Q(csr_gpr_iu_gpr_21__26_) );
	DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_1591_), .Q(csr_gpr_iu_gpr_21__27_) );
	DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_1592_), .Q(csr_gpr_iu_gpr_21__28_) );
	DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_1593_), .Q(csr_gpr_iu_gpr_21__29_) );
	DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_1594_), .Q(csr_gpr_iu_gpr_21__30_) );
	DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_1595_), .Q(csr_gpr_iu_gpr_21__31_) );
	DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_1596_), .Q(csr_gpr_iu_gpr_22__0_) );
	DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_1597_), .Q(csr_gpr_iu_gpr_22__1_) );
	DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_1598_), .Q(csr_gpr_iu_gpr_22__2_) );
	DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_1599_), .Q(csr_gpr_iu_gpr_22__3_) );
	DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_1600_), .Q(csr_gpr_iu_gpr_22__4_) );
	DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_1601_), .Q(csr_gpr_iu_gpr_22__5_) );
	DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_1602_), .Q(csr_gpr_iu_gpr_22__6_) );
	DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_1603_), .Q(csr_gpr_iu_gpr_22__7_) );
	DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_1604_), .Q(csr_gpr_iu_gpr_22__8_) );
	DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_1605_), .Q(csr_gpr_iu_gpr_22__9_) );
	DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_1606_), .Q(csr_gpr_iu_gpr_22__10_) );
	DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_1607_), .Q(csr_gpr_iu_gpr_22__11_) );
	DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_1608_), .Q(csr_gpr_iu_gpr_22__12_) );
	DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_1609_), .Q(csr_gpr_iu_gpr_22__13_) );
	DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_1610_), .Q(csr_gpr_iu_gpr_22__14_) );
	DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_1611_), .Q(csr_gpr_iu_gpr_22__15_) );
	DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_1612_), .Q(csr_gpr_iu_gpr_22__16_) );
	DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_1613_), .Q(csr_gpr_iu_gpr_22__17_) );
	DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_1614_), .Q(csr_gpr_iu_gpr_22__18_) );
	DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_1615_), .Q(csr_gpr_iu_gpr_22__19_) );
	DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_1616_), .Q(csr_gpr_iu_gpr_22__20_) );
	DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_1617_), .Q(csr_gpr_iu_gpr_22__21_) );
	DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_1618_), .Q(csr_gpr_iu_gpr_22__22_) );
	DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_1619_), .Q(csr_gpr_iu_gpr_22__23_) );
	DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_1620_), .Q(csr_gpr_iu_gpr_22__24_) );
	DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_1621_), .Q(csr_gpr_iu_gpr_22__25_) );
	DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_1622_), .Q(csr_gpr_iu_gpr_22__26_) );
	DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_1623_), .Q(csr_gpr_iu_gpr_22__27_) );
	DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_1624_), .Q(csr_gpr_iu_gpr_22__28_) );
	DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_1625_), .Q(csr_gpr_iu_gpr_22__29_) );
	DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_1626_), .Q(csr_gpr_iu_gpr_22__30_) );
	DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1627_), .Q(csr_gpr_iu_gpr_22__31_) );
	DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_2364_), .Q(csr_gpr_iu_gpr_25__0_) );
	DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_2365_), .Q(csr_gpr_iu_gpr_25__1_) );
	DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_2366_), .Q(csr_gpr_iu_gpr_25__2_) );
	DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_2367_), .Q(csr_gpr_iu_gpr_25__3_) );
	DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_2368_), .Q(csr_gpr_iu_gpr_25__4_) );
	DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_2369_), .Q(csr_gpr_iu_gpr_25__5_) );
	DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_2370_), .Q(csr_gpr_iu_gpr_25__6_) );
	DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_2371_), .Q(csr_gpr_iu_gpr_25__7_) );
	DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_2372_), .Q(csr_gpr_iu_gpr_25__8_) );
	DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_2373_), .Q(csr_gpr_iu_gpr_25__9_) );
	DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_2374_), .Q(csr_gpr_iu_gpr_25__10_) );
	DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_2375_), .Q(csr_gpr_iu_gpr_25__11_) );
	DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_2376_), .Q(csr_gpr_iu_gpr_25__12_) );
	DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_2377_), .Q(csr_gpr_iu_gpr_25__13_) );
	DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_2378_), .Q(csr_gpr_iu_gpr_25__14_) );
	DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_2379_), .Q(csr_gpr_iu_gpr_25__15_) );
	DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_2380_), .Q(csr_gpr_iu_gpr_25__16_) );
	DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_2381_), .Q(csr_gpr_iu_gpr_25__17_) );
	DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_2382_), .Q(csr_gpr_iu_gpr_25__18_) );
	DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_2383_), .Q(csr_gpr_iu_gpr_25__19_) );
	DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_2384_), .Q(csr_gpr_iu_gpr_25__20_) );
	DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_2385_), .Q(csr_gpr_iu_gpr_25__21_) );
	DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_2386_), .Q(csr_gpr_iu_gpr_25__22_) );
	DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_2387_), .Q(csr_gpr_iu_gpr_25__23_) );
	DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_2388_), .Q(csr_gpr_iu_gpr_25__24_) );
	DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_2389_), .Q(csr_gpr_iu_gpr_25__25_) );
	DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_2390_), .Q(csr_gpr_iu_gpr_25__26_) );
	DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_2391_), .Q(csr_gpr_iu_gpr_25__27_) );
	DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_2392_), .Q(csr_gpr_iu_gpr_25__28_) );
	DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_2393_), .Q(csr_gpr_iu_gpr_25__29_) );
	DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_2394_), .Q(csr_gpr_iu_gpr_25__30_) );
	DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_2395_), .Q(csr_gpr_iu_gpr_25__31_) );
	DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_1500_), .Q(csr_gpr_iu_gpr_28__0_) );
	DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_1501_), .Q(csr_gpr_iu_gpr_28__1_) );
	DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1502_), .Q(csr_gpr_iu_gpr_28__2_) );
	DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_1503_), .Q(csr_gpr_iu_gpr_28__3_) );
	DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_1504_), .Q(csr_gpr_iu_gpr_28__4_) );
	DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_1505_), .Q(csr_gpr_iu_gpr_28__5_) );
	DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_1506_), .Q(csr_gpr_iu_gpr_28__6_) );
	DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_1507_), .Q(csr_gpr_iu_gpr_28__7_) );
	DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_1508_), .Q(csr_gpr_iu_gpr_28__8_) );
	DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_1509_), .Q(csr_gpr_iu_gpr_28__9_) );
	DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_1510_), .Q(csr_gpr_iu_gpr_28__10_) );
	DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_1511_), .Q(csr_gpr_iu_gpr_28__11_) );
	DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_1512_), .Q(csr_gpr_iu_gpr_28__12_) );
	DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_1513_), .Q(csr_gpr_iu_gpr_28__13_) );
	DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_1514_), .Q(csr_gpr_iu_gpr_28__14_) );
	DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_1515_), .Q(csr_gpr_iu_gpr_28__15_) );
	DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_1516_), .Q(csr_gpr_iu_gpr_28__16_) );
	DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_1517_), .Q(csr_gpr_iu_gpr_28__17_) );
	DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_1518_), .Q(csr_gpr_iu_gpr_28__18_) );
	DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_1519_), .Q(csr_gpr_iu_gpr_28__19_) );
	DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_1520_), .Q(csr_gpr_iu_gpr_28__20_) );
	DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_1521_), .Q(csr_gpr_iu_gpr_28__21_) );
	DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_1522_), .Q(csr_gpr_iu_gpr_28__22_) );
	DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_1523_), .Q(csr_gpr_iu_gpr_28__23_) );
	DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_1524_), .Q(csr_gpr_iu_gpr_28__24_) );
	DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_1525_), .Q(csr_gpr_iu_gpr_28__25_) );
	DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_1526_), .Q(csr_gpr_iu_gpr_28__26_) );
	DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1527_), .Q(csr_gpr_iu_gpr_28__27_) );
	DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_1528_), .Q(csr_gpr_iu_gpr_28__28_) );
	DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_1529_), .Q(csr_gpr_iu_gpr_28__29_) );
	DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_1530_), .Q(csr_gpr_iu_gpr_28__30_) );
	DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_1531_), .Q(csr_gpr_iu_gpr_28__31_) );
	DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_1916_), .Q(csr_gpr_iu_gpr_1__0_) );
	DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_1917_), .Q(csr_gpr_iu_gpr_1__1_) );
	DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1918_), .Q(csr_gpr_iu_gpr_1__2_) );
	DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_1919_), .Q(csr_gpr_iu_gpr_1__3_) );
	DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_1920_), .Q(csr_gpr_iu_gpr_1__4_) );
	DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_1921_), .Q(csr_gpr_iu_gpr_1__5_) );
	DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_1922_), .Q(csr_gpr_iu_gpr_1__6_) );
	DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_1923_), .Q(csr_gpr_iu_gpr_1__7_) );
	DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_1924_), .Q(csr_gpr_iu_gpr_1__8_) );
	DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_1925_), .Q(csr_gpr_iu_gpr_1__9_) );
	DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_1926_), .Q(csr_gpr_iu_gpr_1__10_) );
	DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1927_), .Q(csr_gpr_iu_gpr_1__11_) );
	DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1928_), .Q(csr_gpr_iu_gpr_1__12_) );
	DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1929_), .Q(csr_gpr_iu_gpr_1__13_) );
	DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1930_), .Q(csr_gpr_iu_gpr_1__14_) );
	DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1931_), .Q(csr_gpr_iu_gpr_1__15_) );
	DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1932_), .Q(csr_gpr_iu_gpr_1__16_) );
	DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1933_), .Q(csr_gpr_iu_gpr_1__17_) );
	DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1934_), .Q(csr_gpr_iu_gpr_1__18_) );
	DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1935_), .Q(csr_gpr_iu_gpr_1__19_) );
	DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1936_), .Q(csr_gpr_iu_gpr_1__20_) );
	DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1937_), .Q(csr_gpr_iu_gpr_1__21_) );
	DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1938_), .Q(csr_gpr_iu_gpr_1__22_) );
	DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_1939_), .Q(csr_gpr_iu_gpr_1__23_) );
	DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_1940_), .Q(csr_gpr_iu_gpr_1__24_) );
	DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_1941_), .Q(csr_gpr_iu_gpr_1__25_) );
	DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_1942_), .Q(csr_gpr_iu_gpr_1__26_) );
	DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_1943_), .Q(csr_gpr_iu_gpr_1__27_) );
	DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_1944_), .Q(csr_gpr_iu_gpr_1__28_) );
	DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_1945_), .Q(csr_gpr_iu_gpr_1__29_) );
	DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_1946_), .Q(csr_gpr_iu_gpr_1__30_) );
	DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_1947_), .Q(csr_gpr_iu_gpr_1__31_) );
	DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_1948_), .Q(csr_gpr_iu_gpr_2__0_) );
	DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_1949_), .Q(csr_gpr_iu_gpr_2__1_) );
	DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_1950_), .Q(csr_gpr_iu_gpr_2__2_) );
	DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_1951_), .Q(csr_gpr_iu_gpr_2__3_) );
	DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_1952_), .Q(csr_gpr_iu_gpr_2__4_) );
	DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_1953_), .Q(csr_gpr_iu_gpr_2__5_) );
	DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_1954_), .Q(csr_gpr_iu_gpr_2__6_) );
	DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_1955_), .Q(csr_gpr_iu_gpr_2__7_) );
	DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_1956_), .Q(csr_gpr_iu_gpr_2__8_) );
	DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_1957_), .Q(csr_gpr_iu_gpr_2__9_) );
	DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_1958_), .Q(csr_gpr_iu_gpr_2__10_) );
	DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_1959_), .Q(csr_gpr_iu_gpr_2__11_) );
	DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_1960_), .Q(csr_gpr_iu_gpr_2__12_) );
	DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_1961_), .Q(csr_gpr_iu_gpr_2__13_) );
	DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_1962_), .Q(csr_gpr_iu_gpr_2__14_) );
	DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_1963_), .Q(csr_gpr_iu_gpr_2__15_) );
	DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_1964_), .Q(csr_gpr_iu_gpr_2__16_) );
	DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_1965_), .Q(csr_gpr_iu_gpr_2__17_) );
	DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_1966_), .Q(csr_gpr_iu_gpr_2__18_) );
	DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_1967_), .Q(csr_gpr_iu_gpr_2__19_) );
	DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_1968_), .Q(csr_gpr_iu_gpr_2__20_) );
	DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_1969_), .Q(csr_gpr_iu_gpr_2__21_) );
	DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_1970_), .Q(csr_gpr_iu_gpr_2__22_) );
	DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_1971_), .Q(csr_gpr_iu_gpr_2__23_) );
	DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_1972_), .Q(csr_gpr_iu_gpr_2__24_) );
	DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_1973_), .Q(csr_gpr_iu_gpr_2__25_) );
	DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_1974_), .Q(csr_gpr_iu_gpr_2__26_) );
	DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_1975_), .Q(csr_gpr_iu_gpr_2__27_) );
	DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_1976_), .Q(csr_gpr_iu_gpr_2__28_) );
	DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_1977_), .Q(csr_gpr_iu_gpr_2__29_) );
	DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_1978_), .Q(csr_gpr_iu_gpr_2__30_) );
	DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_1979_), .Q(csr_gpr_iu_gpr_2__31_) );
	DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_1980_), .Q(csr_gpr_iu_gpr_3__0_) );
	DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_1981_), .Q(csr_gpr_iu_gpr_3__1_) );
	DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_1982_), .Q(csr_gpr_iu_gpr_3__2_) );
	DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_1983_), .Q(csr_gpr_iu_gpr_3__3_) );
	DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_1984_), .Q(csr_gpr_iu_gpr_3__4_) );
	DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_1985_), .Q(csr_gpr_iu_gpr_3__5_) );
	DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_1986_), .Q(csr_gpr_iu_gpr_3__6_) );
	DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_1987_), .Q(csr_gpr_iu_gpr_3__7_) );
	DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_1988_), .Q(csr_gpr_iu_gpr_3__8_) );
	DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_1989_), .Q(csr_gpr_iu_gpr_3__9_) );
	DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_1990_), .Q(csr_gpr_iu_gpr_3__10_) );
	DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_1991_), .Q(csr_gpr_iu_gpr_3__11_) );
	DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_1992_), .Q(csr_gpr_iu_gpr_3__12_) );
	DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_1993_), .Q(csr_gpr_iu_gpr_3__13_) );
	DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_1994_), .Q(csr_gpr_iu_gpr_3__14_) );
	DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_1995_), .Q(csr_gpr_iu_gpr_3__15_) );
	DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_1996_), .Q(csr_gpr_iu_gpr_3__16_) );
	DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_1997_), .Q(csr_gpr_iu_gpr_3__17_) );
	DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_1998_), .Q(csr_gpr_iu_gpr_3__18_) );
	DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_1999_), .Q(csr_gpr_iu_gpr_3__19_) );
	DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_2000_), .Q(csr_gpr_iu_gpr_3__20_) );
	DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_2001_), .Q(csr_gpr_iu_gpr_3__21_) );
	DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_2002_), .Q(csr_gpr_iu_gpr_3__22_) );
	DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_2003_), .Q(csr_gpr_iu_gpr_3__23_) );
	DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_2004_), .Q(csr_gpr_iu_gpr_3__24_) );
	DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_2005_), .Q(csr_gpr_iu_gpr_3__25_) );
	DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_2006_), .Q(csr_gpr_iu_gpr_3__26_) );
	DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_2007_), .Q(csr_gpr_iu_gpr_3__27_) );
	DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_2008_), .Q(csr_gpr_iu_gpr_3__28_) );
	DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_2009_), .Q(csr_gpr_iu_gpr_3__29_) );
	DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_2010_), .Q(csr_gpr_iu_gpr_3__30_) );
	DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_2011_), .Q(csr_gpr_iu_gpr_3__31_) );
	DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1756_), .Q(csr_gpr_iu_gpr_14__0_) );
	DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_1757_), .Q(csr_gpr_iu_gpr_14__1_) );
	DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1758_), .Q(csr_gpr_iu_gpr_14__2_) );
	DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1759_), .Q(csr_gpr_iu_gpr_14__3_) );
	DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1760_), .Q(csr_gpr_iu_gpr_14__4_) );
	DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1761_), .Q(csr_gpr_iu_gpr_14__5_) );
	DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1762_), .Q(csr_gpr_iu_gpr_14__6_) );
	DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1763_), .Q(csr_gpr_iu_gpr_14__7_) );
	DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1764_), .Q(csr_gpr_iu_gpr_14__8_) );
	DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1765_), .Q(csr_gpr_iu_gpr_14__9_) );
	DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1766_), .Q(csr_gpr_iu_gpr_14__10_) );
	DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1767_), .Q(csr_gpr_iu_gpr_14__11_) );
	DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1768_), .Q(csr_gpr_iu_gpr_14__12_) );
	DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1769_), .Q(csr_gpr_iu_gpr_14__13_) );
	DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1770_), .Q(csr_gpr_iu_gpr_14__14_) );
	DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1771_), .Q(csr_gpr_iu_gpr_14__15_) );
	DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1772_), .Q(csr_gpr_iu_gpr_14__16_) );
	DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1773_), .Q(csr_gpr_iu_gpr_14__17_) );
	DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1774_), .Q(csr_gpr_iu_gpr_14__18_) );
	DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1775_), .Q(csr_gpr_iu_gpr_14__19_) );
	DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1776_), .Q(csr_gpr_iu_gpr_14__20_) );
	DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1777_), .Q(csr_gpr_iu_gpr_14__21_) );
	DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1778_), .Q(csr_gpr_iu_gpr_14__22_) );
	DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1779_), .Q(csr_gpr_iu_gpr_14__23_) );
	DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1780_), .Q(csr_gpr_iu_gpr_14__24_) );
	DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1781_), .Q(csr_gpr_iu_gpr_14__25_) );
	DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1782_), .Q(csr_gpr_iu_gpr_14__26_) );
	DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1783_), .Q(csr_gpr_iu_gpr_14__27_) );
	DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1784_), .Q(csr_gpr_iu_gpr_14__28_) );
	DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1785_), .Q(csr_gpr_iu_gpr_14__29_) );
	DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1786_), .Q(csr_gpr_iu_gpr_14__30_) );
	DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1787_), .Q(csr_gpr_iu_gpr_14__31_) );
	DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_2012_), .Q(csr_gpr_iu_gpr_4__0_) );
	DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_2013_), .Q(csr_gpr_iu_gpr_4__1_) );
	DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_2014_), .Q(csr_gpr_iu_gpr_4__2_) );
	DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_2015_), .Q(csr_gpr_iu_gpr_4__3_) );
	DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_2016_), .Q(csr_gpr_iu_gpr_4__4_) );
	DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_2017_), .Q(csr_gpr_iu_gpr_4__5_) );
	DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_2018_), .Q(csr_gpr_iu_gpr_4__6_) );
	DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_2019_), .Q(csr_gpr_iu_gpr_4__7_) );
	DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_2020_), .Q(csr_gpr_iu_gpr_4__8_) );
	DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2021_), .Q(csr_gpr_iu_gpr_4__9_) );
	DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_2022_), .Q(csr_gpr_iu_gpr_4__10_) );
	DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_2023_), .Q(csr_gpr_iu_gpr_4__11_) );
	DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_2024_), .Q(csr_gpr_iu_gpr_4__12_) );
	DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_2025_), .Q(csr_gpr_iu_gpr_4__13_) );
	DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2026_), .Q(csr_gpr_iu_gpr_4__14_) );
	DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_2027_), .Q(csr_gpr_iu_gpr_4__15_) );
	DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_2028_), .Q(csr_gpr_iu_gpr_4__16_) );
	DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_2029_), .Q(csr_gpr_iu_gpr_4__17_) );
	DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_2030_), .Q(csr_gpr_iu_gpr_4__18_) );
	DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_2031_), .Q(csr_gpr_iu_gpr_4__19_) );
	DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_2032_), .Q(csr_gpr_iu_gpr_4__20_) );
	DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_2033_), .Q(csr_gpr_iu_gpr_4__21_) );
	DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_2034_), .Q(csr_gpr_iu_gpr_4__22_) );
	DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_2035_), .Q(csr_gpr_iu_gpr_4__23_) );
	DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_2036_), .Q(csr_gpr_iu_gpr_4__24_) );
	DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_2037_), .Q(csr_gpr_iu_gpr_4__25_) );
	DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_2038_), .Q(csr_gpr_iu_gpr_4__26_) );
	DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_2039_), .Q(csr_gpr_iu_gpr_4__27_) );
	DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_2040_), .Q(csr_gpr_iu_gpr_4__28_) );
	DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_2041_), .Q(csr_gpr_iu_gpr_4__29_) );
	DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_2042_), .Q(csr_gpr_iu_gpr_4__30_) );
	DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_2043_), .Q(csr_gpr_iu_gpr_4__31_) );
	DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_2044_), .Q(csr_gpr_iu_gpr_5__0_) );
	DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_2045_), .Q(csr_gpr_iu_gpr_5__1_) );
	DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_2046_), .Q(csr_gpr_iu_gpr_5__2_) );
	DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_2047_), .Q(csr_gpr_iu_gpr_5__3_) );
	DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_2048_), .Q(csr_gpr_iu_gpr_5__4_) );
	DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_2049_), .Q(csr_gpr_iu_gpr_5__5_) );
	DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_2050_), .Q(csr_gpr_iu_gpr_5__6_) );
	DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_2051_), .Q(csr_gpr_iu_gpr_5__7_) );
	DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_2052_), .Q(csr_gpr_iu_gpr_5__8_) );
	DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_2053_), .Q(csr_gpr_iu_gpr_5__9_) );
	DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_2054_), .Q(csr_gpr_iu_gpr_5__10_) );
	DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2055_), .Q(csr_gpr_iu_gpr_5__11_) );
	DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_2056_), .Q(csr_gpr_iu_gpr_5__12_) );
	DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_2057_), .Q(csr_gpr_iu_gpr_5__13_) );
	DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_2058_), .Q(csr_gpr_iu_gpr_5__14_) );
	DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_2059_), .Q(csr_gpr_iu_gpr_5__15_) );
	DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2060_), .Q(csr_gpr_iu_gpr_5__16_) );
	DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2061_), .Q(csr_gpr_iu_gpr_5__17_) );
	DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2062_), .Q(csr_gpr_iu_gpr_5__18_) );
	DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2063_), .Q(csr_gpr_iu_gpr_5__19_) );
	DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2064_), .Q(csr_gpr_iu_gpr_5__20_) );
	DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2065_), .Q(csr_gpr_iu_gpr_5__21_) );
	DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2066_), .Q(csr_gpr_iu_gpr_5__22_) );
	DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2067_), .Q(csr_gpr_iu_gpr_5__23_) );
	DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_2068_), .Q(csr_gpr_iu_gpr_5__24_) );
	DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_2069_), .Q(csr_gpr_iu_gpr_5__25_) );
	DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_2070_), .Q(csr_gpr_iu_gpr_5__26_) );
	DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_2071_), .Q(csr_gpr_iu_gpr_5__27_) );
	DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_2072_), .Q(csr_gpr_iu_gpr_5__28_) );
	DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_2073_), .Q(csr_gpr_iu_gpr_5__29_) );
	DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_2074_), .Q(csr_gpr_iu_gpr_5__30_) );
	DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_2075_), .Q(csr_gpr_iu_gpr_5__31_) );
	DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_2076_), .Q(csr_gpr_iu_gpr_6__0_) );
	DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_2077_), .Q(csr_gpr_iu_gpr_6__1_) );
	DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_2078_), .Q(csr_gpr_iu_gpr_6__2_) );
	DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_2079_), .Q(csr_gpr_iu_gpr_6__3_) );
	DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_2080_), .Q(csr_gpr_iu_gpr_6__4_) );
	DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_2081_), .Q(csr_gpr_iu_gpr_6__5_) );
	DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_2082_), .Q(csr_gpr_iu_gpr_6__6_) );
	DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_2083_), .Q(csr_gpr_iu_gpr_6__7_) );
	DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_2084_), .Q(csr_gpr_iu_gpr_6__8_) );
	DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_2085_), .Q(csr_gpr_iu_gpr_6__9_) );
	DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_2086_), .Q(csr_gpr_iu_gpr_6__10_) );
	DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_2087_), .Q(csr_gpr_iu_gpr_6__11_) );
	DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_2088_), .Q(csr_gpr_iu_gpr_6__12_) );
	DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_2089_), .Q(csr_gpr_iu_gpr_6__13_) );
	DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_2090_), .Q(csr_gpr_iu_gpr_6__14_) );
	DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_2091_), .Q(csr_gpr_iu_gpr_6__15_) );
	DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_2092_), .Q(csr_gpr_iu_gpr_6__16_) );
	DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_2093_), .Q(csr_gpr_iu_gpr_6__17_) );
	DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_2094_), .Q(csr_gpr_iu_gpr_6__18_) );
	DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_2095_), .Q(csr_gpr_iu_gpr_6__19_) );
	DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_2096_), .Q(csr_gpr_iu_gpr_6__20_) );
	DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_2097_), .Q(csr_gpr_iu_gpr_6__21_) );
	DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_2098_), .Q(csr_gpr_iu_gpr_6__22_) );
	DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_2099_), .Q(csr_gpr_iu_gpr_6__23_) );
	DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_2100_), .Q(csr_gpr_iu_gpr_6__24_) );
	DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_2101_), .Q(csr_gpr_iu_gpr_6__25_) );
	DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_2102_), .Q(csr_gpr_iu_gpr_6__26_) );
	DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_2103_), .Q(csr_gpr_iu_gpr_6__27_) );
	DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_2104_), .Q(csr_gpr_iu_gpr_6__28_) );
	DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_2105_), .Q(csr_gpr_iu_gpr_6__29_) );
	DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_2106_), .Q(csr_gpr_iu_gpr_6__30_) );
	DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_2107_), .Q(csr_gpr_iu_gpr_6__31_) );
	DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_2108_), .Q(csr_gpr_iu_gpr_7__0_) );
	DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_2109_), .Q(csr_gpr_iu_gpr_7__1_) );
	DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_2110_), .Q(csr_gpr_iu_gpr_7__2_) );
	DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_2111_), .Q(csr_gpr_iu_gpr_7__3_) );
	DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_2112_), .Q(csr_gpr_iu_gpr_7__4_) );
	DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_2113_), .Q(csr_gpr_iu_gpr_7__5_) );
	DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_2114_), .Q(csr_gpr_iu_gpr_7__6_) );
	DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_2115_), .Q(csr_gpr_iu_gpr_7__7_) );
	DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_2116_), .Q(csr_gpr_iu_gpr_7__8_) );
	DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_2117_), .Q(csr_gpr_iu_gpr_7__9_) );
	DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_2118_), .Q(csr_gpr_iu_gpr_7__10_) );
	DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_2119_), .Q(csr_gpr_iu_gpr_7__11_) );
	DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_2120_), .Q(csr_gpr_iu_gpr_7__12_) );
	DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_2121_), .Q(csr_gpr_iu_gpr_7__13_) );
	DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_2122_), .Q(csr_gpr_iu_gpr_7__14_) );
	DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_2123_), .Q(csr_gpr_iu_gpr_7__15_) );
	DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_2124_), .Q(csr_gpr_iu_gpr_7__16_) );
	DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_2125_), .Q(csr_gpr_iu_gpr_7__17_) );
	DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_2126_), .Q(csr_gpr_iu_gpr_7__18_) );
	DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_2127_), .Q(csr_gpr_iu_gpr_7__19_) );
	DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_2128_), .Q(csr_gpr_iu_gpr_7__20_) );
	DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_2129_), .Q(csr_gpr_iu_gpr_7__21_) );
	DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_2130_), .Q(csr_gpr_iu_gpr_7__22_) );
	DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_2131_), .Q(csr_gpr_iu_gpr_7__23_) );
	DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_2132_), .Q(csr_gpr_iu_gpr_7__24_) );
	DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_2133_), .Q(csr_gpr_iu_gpr_7__25_) );
	DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_2134_), .Q(csr_gpr_iu_gpr_7__26_) );
	DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_2135_), .Q(csr_gpr_iu_gpr_7__27_) );
	DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_2136_), .Q(csr_gpr_iu_gpr_7__28_) );
	DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_2137_), .Q(csr_gpr_iu_gpr_7__29_) );
	DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_2138_), .Q(csr_gpr_iu_gpr_7__30_) );
	DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_2139_), .Q(csr_gpr_iu_gpr_7__31_) );
	DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_1820_), .Q(csr_gpr_iu_gpr_15__0_) );
	DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1821_), .Q(csr_gpr_iu_gpr_15__1_) );
	DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_1822_), .Q(csr_gpr_iu_gpr_15__2_) );
	DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1823_), .Q(csr_gpr_iu_gpr_15__3_) );
	DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1824_), .Q(csr_gpr_iu_gpr_15__4_) );
	DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1825_), .Q(csr_gpr_iu_gpr_15__5_) );
	DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1826_), .Q(csr_gpr_iu_gpr_15__6_) );
	DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1827_), .Q(csr_gpr_iu_gpr_15__7_) );
	DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1828_), .Q(csr_gpr_iu_gpr_15__8_) );
	DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1829_), .Q(csr_gpr_iu_gpr_15__9_) );
	DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1830_), .Q(csr_gpr_iu_gpr_15__10_) );
	DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1831_), .Q(csr_gpr_iu_gpr_15__11_) );
	DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1832_), .Q(csr_gpr_iu_gpr_15__12_) );
	DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1833_), .Q(csr_gpr_iu_gpr_15__13_) );
	DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1834_), .Q(csr_gpr_iu_gpr_15__14_) );
	DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1835_), .Q(csr_gpr_iu_gpr_15__15_) );
	DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1836_), .Q(csr_gpr_iu_gpr_15__16_) );
	DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1837_), .Q(csr_gpr_iu_gpr_15__17_) );
	DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1838_), .Q(csr_gpr_iu_gpr_15__18_) );
	DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1839_), .Q(csr_gpr_iu_gpr_15__19_) );
	DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1840_), .Q(csr_gpr_iu_gpr_15__20_) );
	DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1841_), .Q(csr_gpr_iu_gpr_15__21_) );
	DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1842_), .Q(csr_gpr_iu_gpr_15__22_) );
	DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1843_), .Q(csr_gpr_iu_gpr_15__23_) );
	DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1844_), .Q(csr_gpr_iu_gpr_15__24_) );
	DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1845_), .Q(csr_gpr_iu_gpr_15__25_) );
	DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1846_), .Q(csr_gpr_iu_gpr_15__26_) );
	DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1847_), .Q(csr_gpr_iu_gpr_15__27_) );
	DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1848_), .Q(csr_gpr_iu_gpr_15__28_) );
	DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1849_), .Q(csr_gpr_iu_gpr_15__29_) );
	DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1850_), .Q(csr_gpr_iu_gpr_15__30_) );
	DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1851_), .Q(csr_gpr_iu_gpr_15__31_) );
	DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_2140_), .Q(csr_gpr_iu_gpr_8__0_) );
	DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_2141_), .Q(csr_gpr_iu_gpr_8__1_) );
	DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_2142_), .Q(csr_gpr_iu_gpr_8__2_) );
	DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_2143_), .Q(csr_gpr_iu_gpr_8__3_) );
	DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_2144_), .Q(csr_gpr_iu_gpr_8__4_) );
	DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_2145_), .Q(csr_gpr_iu_gpr_8__5_) );
	DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_2146_), .Q(csr_gpr_iu_gpr_8__6_) );
	DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_2147_), .Q(csr_gpr_iu_gpr_8__7_) );
	DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_2148_), .Q(csr_gpr_iu_gpr_8__8_) );
	DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_2149_), .Q(csr_gpr_iu_gpr_8__9_) );
	DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2150_), .Q(csr_gpr_iu_gpr_8__10_) );
	DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_2151_), .Q(csr_gpr_iu_gpr_8__11_) );
	DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_2152_), .Q(csr_gpr_iu_gpr_8__12_) );
	DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_2153_), .Q(csr_gpr_iu_gpr_8__13_) );
	DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_2154_), .Q(csr_gpr_iu_gpr_8__14_) );
	DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2155_), .Q(csr_gpr_iu_gpr_8__15_) );
	DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_2156_), .Q(csr_gpr_iu_gpr_8__16_) );
	DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_2157_), .Q(csr_gpr_iu_gpr_8__17_) );
	DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_2158_), .Q(csr_gpr_iu_gpr_8__18_) );
	DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_2159_), .Q(csr_gpr_iu_gpr_8__19_) );
	DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_2160_), .Q(csr_gpr_iu_gpr_8__20_) );
	DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_2161_), .Q(csr_gpr_iu_gpr_8__21_) );
	DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_2162_), .Q(csr_gpr_iu_gpr_8__22_) );
	DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_2163_), .Q(csr_gpr_iu_gpr_8__23_) );
	DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_2164_), .Q(csr_gpr_iu_gpr_8__24_) );
	DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_2165_), .Q(csr_gpr_iu_gpr_8__25_) );
	DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_2166_), .Q(csr_gpr_iu_gpr_8__26_) );
	DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_2167_), .Q(csr_gpr_iu_gpr_8__27_) );
	DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_2168_), .Q(csr_gpr_iu_gpr_8__28_) );
	DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_2169_), .Q(csr_gpr_iu_gpr_8__29_) );
	DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_2170_), .Q(csr_gpr_iu_gpr_8__30_) );
	DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_2171_), .Q(csr_gpr_iu_gpr_8__31_) );
	DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_2236_), .Q(csr_gpr_iu_gpr_9__0_) );
	DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_2237_), .Q(csr_gpr_iu_gpr_9__1_) );
	DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_2238_), .Q(csr_gpr_iu_gpr_9__2_) );
	DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_2239_), .Q(csr_gpr_iu_gpr_9__3_) );
	DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_2240_), .Q(csr_gpr_iu_gpr_9__4_) );
	DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_2241_), .Q(csr_gpr_iu_gpr_9__5_) );
	DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_2242_), .Q(csr_gpr_iu_gpr_9__6_) );
	DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_2243_), .Q(csr_gpr_iu_gpr_9__7_) );
	DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_2244_), .Q(csr_gpr_iu_gpr_9__8_) );
	DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_2245_), .Q(csr_gpr_iu_gpr_9__9_) );
	DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_2246_), .Q(csr_gpr_iu_gpr_9__10_) );
	DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_2247_), .Q(csr_gpr_iu_gpr_9__11_) );
	DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_2248_), .Q(csr_gpr_iu_gpr_9__12_) );
	DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_2249_), .Q(csr_gpr_iu_gpr_9__13_) );
	DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_2250_), .Q(csr_gpr_iu_gpr_9__14_) );
	DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_2251_), .Q(csr_gpr_iu_gpr_9__15_) );
	DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_2252_), .Q(csr_gpr_iu_gpr_9__16_) );
	DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2253_), .Q(csr_gpr_iu_gpr_9__17_) );
	DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2254_), .Q(csr_gpr_iu_gpr_9__18_) );
	DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2255_), .Q(csr_gpr_iu_gpr_9__19_) );
	DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2256_), .Q(csr_gpr_iu_gpr_9__20_) );
	DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2257_), .Q(csr_gpr_iu_gpr_9__21_) );
	DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2258_), .Q(csr_gpr_iu_gpr_9__22_) );
	DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2259_), .Q(csr_gpr_iu_gpr_9__23_) );
	DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2260_), .Q(csr_gpr_iu_gpr_9__24_) );
	DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_2261_), .Q(csr_gpr_iu_gpr_9__25_) );
	DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_2262_), .Q(csr_gpr_iu_gpr_9__26_) );
	DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_2263_), .Q(csr_gpr_iu_gpr_9__27_) );
	DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_2264_), .Q(csr_gpr_iu_gpr_9__28_) );
	DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_2265_), .Q(csr_gpr_iu_gpr_9__29_) );
	DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_2266_), .Q(csr_gpr_iu_gpr_9__30_) );
	DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_2267_), .Q(csr_gpr_iu_gpr_9__31_) );
	DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_2268_), .Q(csr_gpr_iu_gpr_10__0_) );
	DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_2269_), .Q(csr_gpr_iu_gpr_10__1_) );
	DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_2270_), .Q(csr_gpr_iu_gpr_10__2_) );
	DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_2271_), .Q(csr_gpr_iu_gpr_10__3_) );
	DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_2272_), .Q(csr_gpr_iu_gpr_10__4_) );
	DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_2273_), .Q(csr_gpr_iu_gpr_10__5_) );
	DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_2274_), .Q(csr_gpr_iu_gpr_10__6_) );
	DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_2275_), .Q(csr_gpr_iu_gpr_10__7_) );
	DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_2276_), .Q(csr_gpr_iu_gpr_10__8_) );
	DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_2277_), .Q(csr_gpr_iu_gpr_10__9_) );
	DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_2278_), .Q(csr_gpr_iu_gpr_10__10_) );
	DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_2279_), .Q(csr_gpr_iu_gpr_10__11_) );
	DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_2280_), .Q(csr_gpr_iu_gpr_10__12_) );
	DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_2281_), .Q(csr_gpr_iu_gpr_10__13_) );
	DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_2282_), .Q(csr_gpr_iu_gpr_10__14_) );
	DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_2283_), .Q(csr_gpr_iu_gpr_10__15_) );
	DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_2284_), .Q(csr_gpr_iu_gpr_10__16_) );
	DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_2285_), .Q(csr_gpr_iu_gpr_10__17_) );
	DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_2286_), .Q(csr_gpr_iu_gpr_10__18_) );
	DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_2287_), .Q(csr_gpr_iu_gpr_10__19_) );
	DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_2288_), .Q(csr_gpr_iu_gpr_10__20_) );
	DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_2289_), .Q(csr_gpr_iu_gpr_10__21_) );
	DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_2290_), .Q(csr_gpr_iu_gpr_10__22_) );
	DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_2291_), .Q(csr_gpr_iu_gpr_10__23_) );
	DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_2292_), .Q(csr_gpr_iu_gpr_10__24_) );
	DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_2293_), .Q(csr_gpr_iu_gpr_10__25_) );
	DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_2294_), .Q(csr_gpr_iu_gpr_10__26_) );
	DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_2295_), .Q(csr_gpr_iu_gpr_10__27_) );
	DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_2296_), .Q(csr_gpr_iu_gpr_10__28_) );
	DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_2297_), .Q(csr_gpr_iu_gpr_10__29_) );
	DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_2298_), .Q(csr_gpr_iu_gpr_10__30_) );
	DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_2299_), .Q(csr_gpr_iu_gpr_10__31_) );
	DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_2300_), .Q(csr_gpr_iu_gpr_11__0_) );
	DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_2301_), .Q(csr_gpr_iu_gpr_11__1_) );
	DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_2302_), .Q(csr_gpr_iu_gpr_11__2_) );
	DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_2303_), .Q(csr_gpr_iu_gpr_11__3_) );
	DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_2304_), .Q(csr_gpr_iu_gpr_11__4_) );
	DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_2305_), .Q(csr_gpr_iu_gpr_11__5_) );
	DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_2306_), .Q(csr_gpr_iu_gpr_11__6_) );
	DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_2307_), .Q(csr_gpr_iu_gpr_11__7_) );
	DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_2308_), .Q(csr_gpr_iu_gpr_11__8_) );
	DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_2309_), .Q(csr_gpr_iu_gpr_11__9_) );
	DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_2310_), .Q(csr_gpr_iu_gpr_11__10_) );
	DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_2311_), .Q(csr_gpr_iu_gpr_11__11_) );
	DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_2312_), .Q(csr_gpr_iu_gpr_11__12_) );
	DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_2313_), .Q(csr_gpr_iu_gpr_11__13_) );
	DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_2314_), .Q(csr_gpr_iu_gpr_11__14_) );
	DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_2315_), .Q(csr_gpr_iu_gpr_11__15_) );
	DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_2316_), .Q(csr_gpr_iu_gpr_11__16_) );
	DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_2317_), .Q(csr_gpr_iu_gpr_11__17_) );
	DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_2318_), .Q(csr_gpr_iu_gpr_11__18_) );
	DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_2319_), .Q(csr_gpr_iu_gpr_11__19_) );
	DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_2320_), .Q(csr_gpr_iu_gpr_11__20_) );
	DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_2321_), .Q(csr_gpr_iu_gpr_11__21_) );
	DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_2322_), .Q(csr_gpr_iu_gpr_11__22_) );
	DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_2323_), .Q(csr_gpr_iu_gpr_11__23_) );
	DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_2324_), .Q(csr_gpr_iu_gpr_11__24_) );
	DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_2325_), .Q(csr_gpr_iu_gpr_11__25_) );
	DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_2326_), .Q(csr_gpr_iu_gpr_11__26_) );
	DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_2327_), .Q(csr_gpr_iu_gpr_11__27_) );
	DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_2328_), .Q(csr_gpr_iu_gpr_11__28_) );
	DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_2329_), .Q(csr_gpr_iu_gpr_11__29_) );
	DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_2330_), .Q(csr_gpr_iu_gpr_11__30_) );
	DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_2331_), .Q(csr_gpr_iu_gpr_11__31_) );
	DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_1884_), .Q(csr_gpr_iu_gpr_0__0_) );
	DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_1885_), .Q(csr_gpr_iu_gpr_0__1_) );
	DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1886_), .Q(csr_gpr_iu_gpr_0__2_) );
	DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_1887_), .Q(csr_gpr_iu_gpr_0__3_) );
	DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1888_), .Q(csr_gpr_iu_gpr_0__4_) );
	DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1889_), .Q(csr_gpr_iu_gpr_0__5_) );
	DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1890_), .Q(csr_gpr_iu_gpr_0__6_) );
	DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1891_), .Q(csr_gpr_iu_gpr_0__7_) );
	DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1892_), .Q(csr_gpr_iu_gpr_0__8_) );
	DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1893_), .Q(csr_gpr_iu_gpr_0__9_) );
	DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1894_), .Q(csr_gpr_iu_gpr_0__10_) );
	DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1895_), .Q(csr_gpr_iu_gpr_0__11_) );
	DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1896_), .Q(csr_gpr_iu_gpr_0__12_) );
	DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1897_), .Q(csr_gpr_iu_gpr_0__13_) );
	DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1898_), .Q(csr_gpr_iu_gpr_0__14_) );
	DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1899_), .Q(csr_gpr_iu_gpr_0__15_) );
	DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1900_), .Q(csr_gpr_iu_gpr_0__16_) );
	DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1901_), .Q(csr_gpr_iu_gpr_0__17_) );
	DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1902_), .Q(csr_gpr_iu_gpr_0__18_) );
	DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1903_), .Q(csr_gpr_iu_gpr_0__19_) );
	DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1904_), .Q(csr_gpr_iu_gpr_0__20_) );
	DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1905_), .Q(csr_gpr_iu_gpr_0__21_) );
	DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1906_), .Q(csr_gpr_iu_gpr_0__22_) );
	DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1907_), .Q(csr_gpr_iu_gpr_0__23_) );
	DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1908_), .Q(csr_gpr_iu_gpr_0__24_) );
	DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1909_), .Q(csr_gpr_iu_gpr_0__25_) );
	DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1910_), .Q(csr_gpr_iu_gpr_0__26_) );
	DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1911_), .Q(csr_gpr_iu_gpr_0__27_) );
	DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1912_), .Q(csr_gpr_iu_gpr_0__28_) );
	DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1913_), .Q(csr_gpr_iu_gpr_0__29_) );
	DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1914_), .Q(csr_gpr_iu_gpr_0__30_) );
	DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1915_), .Q(csr_gpr_iu_gpr_0__31_) );
	DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_2172_), .Q(csr_gpr_iu_gpr_12__0_) );
	DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_2173_), .Q(csr_gpr_iu_gpr_12__1_) );
	DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_2174_), .Q(csr_gpr_iu_gpr_12__2_) );
	DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_2175_), .Q(csr_gpr_iu_gpr_12__3_) );
	DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_2176_), .Q(csr_gpr_iu_gpr_12__4_) );
	DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_2177_), .Q(csr_gpr_iu_gpr_12__5_) );
	DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_2178_), .Q(csr_gpr_iu_gpr_12__6_) );
	DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_2179_), .Q(csr_gpr_iu_gpr_12__7_) );
	DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_2180_), .Q(csr_gpr_iu_gpr_12__8_) );
	DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_2181_), .Q(csr_gpr_iu_gpr_12__9_) );
	DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_2182_), .Q(csr_gpr_iu_gpr_12__10_) );
	DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2183_), .Q(csr_gpr_iu_gpr_12__11_) );
	DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_2184_), .Q(csr_gpr_iu_gpr_12__12_) );
	DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_2185_), .Q(csr_gpr_iu_gpr_12__13_) );
	DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_2186_), .Q(csr_gpr_iu_gpr_12__14_) );
	DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_2187_), .Q(csr_gpr_iu_gpr_12__15_) );
	DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2188_), .Q(csr_gpr_iu_gpr_12__16_) );
	DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_2189_), .Q(csr_gpr_iu_gpr_12__17_) );
	DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_2190_), .Q(csr_gpr_iu_gpr_12__18_) );
	DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_2191_), .Q(csr_gpr_iu_gpr_12__19_) );
	DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_2192_), .Q(csr_gpr_iu_gpr_12__20_) );
	DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_2193_), .Q(csr_gpr_iu_gpr_12__21_) );
	DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_2194_), .Q(csr_gpr_iu_gpr_12__22_) );
	DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_2195_), .Q(csr_gpr_iu_gpr_12__23_) );
	DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_2196_), .Q(csr_gpr_iu_gpr_12__24_) );
	DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_2197_), .Q(csr_gpr_iu_gpr_12__25_) );
	DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_2198_), .Q(csr_gpr_iu_gpr_12__26_) );
	DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_2199_), .Q(csr_gpr_iu_gpr_12__27_) );
	DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_2200_), .Q(csr_gpr_iu_gpr_12__28_) );
	DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_2201_), .Q(csr_gpr_iu_gpr_12__29_) );
	DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_2202_), .Q(csr_gpr_iu_gpr_12__30_) );
	DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_2203_), .Q(csr_gpr_iu_gpr_12__31_) );
	DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_1724_), .Q(csr_gpr_iu_gpr_19__0_) );
	DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_1725_), .Q(csr_gpr_iu_gpr_19__1_) );
	DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_1726_), .Q(csr_gpr_iu_gpr_19__2_) );
	DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_1727_), .Q(csr_gpr_iu_gpr_19__3_) );
	DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_1728_), .Q(csr_gpr_iu_gpr_19__4_) );
	DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1729_), .Q(csr_gpr_iu_gpr_19__5_) );
	DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_1730_), .Q(csr_gpr_iu_gpr_19__6_) );
	DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_1731_), .Q(csr_gpr_iu_gpr_19__7_) );
	DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_1732_), .Q(csr_gpr_iu_gpr_19__8_) );
	DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_1733_), .Q(csr_gpr_iu_gpr_19__9_) );
	DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_1734_), .Q(csr_gpr_iu_gpr_19__10_) );
	DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_1735_), .Q(csr_gpr_iu_gpr_19__11_) );
	DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_1736_), .Q(csr_gpr_iu_gpr_19__12_) );
	DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_1737_), .Q(csr_gpr_iu_gpr_19__13_) );
	DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1738_), .Q(csr_gpr_iu_gpr_19__14_) );
	DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1739_), .Q(csr_gpr_iu_gpr_19__15_) );
	DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1740_), .Q(csr_gpr_iu_gpr_19__16_) );
	DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1741_), .Q(csr_gpr_iu_gpr_19__17_) );
	DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1742_), .Q(csr_gpr_iu_gpr_19__18_) );
	DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1743_), .Q(csr_gpr_iu_gpr_19__19_) );
	DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1744_), .Q(csr_gpr_iu_gpr_19__20_) );
	DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1745_), .Q(csr_gpr_iu_gpr_19__21_) );
	DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1746_), .Q(csr_gpr_iu_gpr_19__22_) );
	DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1747_), .Q(csr_gpr_iu_gpr_19__23_) );
	DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1748_), .Q(csr_gpr_iu_gpr_19__24_) );
	DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1749_), .Q(csr_gpr_iu_gpr_19__25_) );
	DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_1750_), .Q(csr_gpr_iu_gpr_19__26_) );
	DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_1751_), .Q(csr_gpr_iu_gpr_19__27_) );
	DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_1752_), .Q(csr_gpr_iu_gpr_19__28_) );
	DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_1753_), .Q(csr_gpr_iu_gpr_19__29_) );
	DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_1754_), .Q(csr_gpr_iu_gpr_19__30_) );
	DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_1755_), .Q(csr_gpr_iu_gpr_19__31_) );
	DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_1788_), .Q(csr_gpr_iu_gpr_16__0_) );
	DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_1789_), .Q(csr_gpr_iu_gpr_16__1_) );
	DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_1790_), .Q(csr_gpr_iu_gpr_16__2_) );
	DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_1791_), .Q(csr_gpr_iu_gpr_16__3_) );
	DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_1792_), .Q(csr_gpr_iu_gpr_16__4_) );
	DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_1793_), .Q(csr_gpr_iu_gpr_16__5_) );
	DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_1794_), .Q(csr_gpr_iu_gpr_16__6_) );
	DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_1795_), .Q(csr_gpr_iu_gpr_16__7_) );
	DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_1796_), .Q(csr_gpr_iu_gpr_16__8_) );
	DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_1797_), .Q(csr_gpr_iu_gpr_16__9_) );
	DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_1798_), .Q(csr_gpr_iu_gpr_16__10_) );
	DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_1799_), .Q(csr_gpr_iu_gpr_16__11_) );
	DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_1800_), .Q(csr_gpr_iu_gpr_16__12_) );
	DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_1801_), .Q(csr_gpr_iu_gpr_16__13_) );
	DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_1802_), .Q(csr_gpr_iu_gpr_16__14_) );
	DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_1803_), .Q(csr_gpr_iu_gpr_16__15_) );
	DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_1804_), .Q(csr_gpr_iu_gpr_16__16_) );
	DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_1805_), .Q(csr_gpr_iu_gpr_16__17_) );
	DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_1806_), .Q(csr_gpr_iu_gpr_16__18_) );
	DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_1807_), .Q(csr_gpr_iu_gpr_16__19_) );
	DFFPOSX1 DFFPOSX1_993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_1808_), .Q(csr_gpr_iu_gpr_16__20_) );
	DFFPOSX1 DFFPOSX1_994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_1809_), .Q(csr_gpr_iu_gpr_16__21_) );
	DFFPOSX1 DFFPOSX1_995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_1810_), .Q(csr_gpr_iu_gpr_16__22_) );
	DFFPOSX1 DFFPOSX1_996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_1811_), .Q(csr_gpr_iu_gpr_16__23_) );
	DFFPOSX1 DFFPOSX1_997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_1812_), .Q(csr_gpr_iu_gpr_16__24_) );
	DFFPOSX1 DFFPOSX1_998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_1813_), .Q(csr_gpr_iu_gpr_16__25_) );
	DFFPOSX1 DFFPOSX1_999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_1814_), .Q(csr_gpr_iu_gpr_16__26_) );
	DFFPOSX1 DFFPOSX1_1000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_1815_), .Q(csr_gpr_iu_gpr_16__27_) );
	DFFPOSX1 DFFPOSX1_1001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_1816_), .Q(csr_gpr_iu_gpr_16__28_) );
	DFFPOSX1 DFFPOSX1_1002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_1817_), .Q(csr_gpr_iu_gpr_16__29_) );
	DFFPOSX1 DFFPOSX1_1003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_1818_), .Q(csr_gpr_iu_gpr_16__30_) );
	DFFPOSX1 DFFPOSX1_1004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_1819_), .Q(csr_gpr_iu_gpr_16__31_) );
	DFFPOSX1 DFFPOSX1_1005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_1852_), .Q(csr_gpr_iu_gpr_17__0_) );
	DFFPOSX1 DFFPOSX1_1006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_1853_), .Q(csr_gpr_iu_gpr_17__1_) );
	DFFPOSX1 DFFPOSX1_1007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_1854_), .Q(csr_gpr_iu_gpr_17__2_) );
	DFFPOSX1 DFFPOSX1_1008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_1855_), .Q(csr_gpr_iu_gpr_17__3_) );
	DFFPOSX1 DFFPOSX1_1009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_1856_), .Q(csr_gpr_iu_gpr_17__4_) );
	DFFPOSX1 DFFPOSX1_1010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_1857_), .Q(csr_gpr_iu_gpr_17__5_) );
	DFFPOSX1 DFFPOSX1_1011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_1858_), .Q(csr_gpr_iu_gpr_17__6_) );
	DFFPOSX1 DFFPOSX1_1012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_1859_), .Q(csr_gpr_iu_gpr_17__7_) );
	DFFPOSX1 DFFPOSX1_1013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_1860_), .Q(csr_gpr_iu_gpr_17__8_) );
	DFFPOSX1 DFFPOSX1_1014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_1861_), .Q(csr_gpr_iu_gpr_17__9_) );
	DFFPOSX1 DFFPOSX1_1015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_1862_), .Q(csr_gpr_iu_gpr_17__10_) );
	DFFPOSX1 DFFPOSX1_1016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_1863_), .Q(csr_gpr_iu_gpr_17__11_) );
	DFFPOSX1 DFFPOSX1_1017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_1864_), .Q(csr_gpr_iu_gpr_17__12_) );
	DFFPOSX1 DFFPOSX1_1018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_1865_), .Q(csr_gpr_iu_gpr_17__13_) );
	DFFPOSX1 DFFPOSX1_1019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_1866_), .Q(csr_gpr_iu_gpr_17__14_) );
	DFFPOSX1 DFFPOSX1_1020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_1867_), .Q(csr_gpr_iu_gpr_17__15_) );
	DFFPOSX1 DFFPOSX1_1021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_1868_), .Q(csr_gpr_iu_gpr_17__16_) );
	DFFPOSX1 DFFPOSX1_1022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_1869_), .Q(csr_gpr_iu_gpr_17__17_) );
	DFFPOSX1 DFFPOSX1_1023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_1870_), .Q(csr_gpr_iu_gpr_17__18_) );
	DFFPOSX1 DFFPOSX1_1024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_1871_), .Q(csr_gpr_iu_gpr_17__19_) );
	DFFPOSX1 DFFPOSX1_1025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_1872_), .Q(csr_gpr_iu_gpr_17__20_) );
	DFFPOSX1 DFFPOSX1_1026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_1873_), .Q(csr_gpr_iu_gpr_17__21_) );
	DFFPOSX1 DFFPOSX1_1027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_1874_), .Q(csr_gpr_iu_gpr_17__22_) );
	DFFPOSX1 DFFPOSX1_1028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_1875_), .Q(csr_gpr_iu_gpr_17__23_) );
	DFFPOSX1 DFFPOSX1_1029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_1876_), .Q(csr_gpr_iu_gpr_17__24_) );
	DFFPOSX1 DFFPOSX1_1030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_1877_), .Q(csr_gpr_iu_gpr_17__25_) );
	DFFPOSX1 DFFPOSX1_1031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_1878_), .Q(csr_gpr_iu_gpr_17__26_) );
	DFFPOSX1 DFFPOSX1_1032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_1879_), .Q(csr_gpr_iu_gpr_17__27_) );
	DFFPOSX1 DFFPOSX1_1033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_1880_), .Q(csr_gpr_iu_gpr_17__28_) );
	DFFPOSX1 DFFPOSX1_1034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_1881_), .Q(csr_gpr_iu_gpr_17__29_) );
	DFFPOSX1 DFFPOSX1_1035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_1882_), .Q(csr_gpr_iu_gpr_17__30_) );
	DFFPOSX1 DFFPOSX1_1036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_1883_), .Q(csr_gpr_iu_gpr_17__31_) );
	DFFPOSX1 DFFPOSX1_1037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_1468_), .Q(csr_gpr_iu_gpr_30__0_) );
	DFFPOSX1 DFFPOSX1_1038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_1469_), .Q(csr_gpr_iu_gpr_30__1_) );
	DFFPOSX1 DFFPOSX1_1039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_1470_), .Q(csr_gpr_iu_gpr_30__2_) );
	DFFPOSX1 DFFPOSX1_1040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_1471_), .Q(csr_gpr_iu_gpr_30__3_) );
	DFFPOSX1 DFFPOSX1_1041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_1472_), .Q(csr_gpr_iu_gpr_30__4_) );
	DFFPOSX1 DFFPOSX1_1042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1473_), .Q(csr_gpr_iu_gpr_30__5_) );
	DFFPOSX1 DFFPOSX1_1043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1474_), .Q(csr_gpr_iu_gpr_30__6_) );
	DFFPOSX1 DFFPOSX1_1044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1475_), .Q(csr_gpr_iu_gpr_30__7_) );
	DFFPOSX1 DFFPOSX1_1045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1476_), .Q(csr_gpr_iu_gpr_30__8_) );
	DFFPOSX1 DFFPOSX1_1046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1477_), .Q(csr_gpr_iu_gpr_30__9_) );
	DFFPOSX1 DFFPOSX1_1047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1478_), .Q(csr_gpr_iu_gpr_30__10_) );
	DFFPOSX1 DFFPOSX1_1048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1479_), .Q(csr_gpr_iu_gpr_30__11_) );
	DFFPOSX1 DFFPOSX1_1049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1480_), .Q(csr_gpr_iu_gpr_30__12_) );
	DFFPOSX1 DFFPOSX1_1050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1481_), .Q(csr_gpr_iu_gpr_30__13_) );
	DFFPOSX1 DFFPOSX1_1051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1482_), .Q(csr_gpr_iu_gpr_30__14_) );
	DFFPOSX1 DFFPOSX1_1052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1483_), .Q(csr_gpr_iu_gpr_30__15_) );
	DFFPOSX1 DFFPOSX1_1053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1484_), .Q(csr_gpr_iu_gpr_30__16_) );
	DFFPOSX1 DFFPOSX1_1054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1485_), .Q(csr_gpr_iu_gpr_30__17_) );
	DFFPOSX1 DFFPOSX1_1055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1486_), .Q(csr_gpr_iu_gpr_30__18_) );
	DFFPOSX1 DFFPOSX1_1056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1487_), .Q(csr_gpr_iu_gpr_30__19_) );
	DFFPOSX1 DFFPOSX1_1057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1488_), .Q(csr_gpr_iu_gpr_30__20_) );
	DFFPOSX1 DFFPOSX1_1058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1489_), .Q(csr_gpr_iu_gpr_30__21_) );
	DFFPOSX1 DFFPOSX1_1059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1490_), .Q(csr_gpr_iu_gpr_30__22_) );
	DFFPOSX1 DFFPOSX1_1060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1491_), .Q(csr_gpr_iu_gpr_30__23_) );
	DFFPOSX1 DFFPOSX1_1061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1492_), .Q(csr_gpr_iu_gpr_30__24_) );
	DFFPOSX1 DFFPOSX1_1062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1493_), .Q(csr_gpr_iu_gpr_30__25_) );
	DFFPOSX1 DFFPOSX1_1063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1494_), .Q(csr_gpr_iu_gpr_30__26_) );
	DFFPOSX1 DFFPOSX1_1064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1495_), .Q(csr_gpr_iu_gpr_30__27_) );
	DFFPOSX1 DFFPOSX1_1065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1496_), .Q(csr_gpr_iu_gpr_30__28_) );
	DFFPOSX1 DFFPOSX1_1066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1497_), .Q(csr_gpr_iu_gpr_30__29_) );
	DFFPOSX1 DFFPOSX1_1067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1498_), .Q(csr_gpr_iu_gpr_30__30_) );
	DFFPOSX1 DFFPOSX1_1068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1499_), .Q(csr_gpr_iu_gpr_30__31_) );
	DFFPOSX1 DFFPOSX1_1069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1660_), .Q(csr_gpr_iu_gpr_24__0_) );
	DFFPOSX1 DFFPOSX1_1070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1661_), .Q(csr_gpr_iu_gpr_24__1_) );
	DFFPOSX1 DFFPOSX1_1071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1662_), .Q(csr_gpr_iu_gpr_24__2_) );
	DFFPOSX1 DFFPOSX1_1072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_1663_), .Q(csr_gpr_iu_gpr_24__3_) );
	DFFPOSX1 DFFPOSX1_1073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_1664_), .Q(csr_gpr_iu_gpr_24__4_) );
	DFFPOSX1 DFFPOSX1_1074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_1665_), .Q(csr_gpr_iu_gpr_24__5_) );
	DFFPOSX1 DFFPOSX1_1075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_1666_), .Q(csr_gpr_iu_gpr_24__6_) );
	DFFPOSX1 DFFPOSX1_1076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_1667_), .Q(csr_gpr_iu_gpr_24__7_) );
	DFFPOSX1 DFFPOSX1_1077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_1668_), .Q(csr_gpr_iu_gpr_24__8_) );
	DFFPOSX1 DFFPOSX1_1078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_1669_), .Q(csr_gpr_iu_gpr_24__9_) );
	DFFPOSX1 DFFPOSX1_1079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_1670_), .Q(csr_gpr_iu_gpr_24__10_) );
	DFFPOSX1 DFFPOSX1_1080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_1671_), .Q(csr_gpr_iu_gpr_24__11_) );
	DFFPOSX1 DFFPOSX1_1081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_1672_), .Q(csr_gpr_iu_gpr_24__12_) );
	DFFPOSX1 DFFPOSX1_1082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_1673_), .Q(csr_gpr_iu_gpr_24__13_) );
	DFFPOSX1 DFFPOSX1_1083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_1674_), .Q(csr_gpr_iu_gpr_24__14_) );
	DFFPOSX1 DFFPOSX1_1084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_1675_), .Q(csr_gpr_iu_gpr_24__15_) );
	DFFPOSX1 DFFPOSX1_1085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_1676_), .Q(csr_gpr_iu_gpr_24__16_) );
	DFFPOSX1 DFFPOSX1_1086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_1677_), .Q(csr_gpr_iu_gpr_24__17_) );
	DFFPOSX1 DFFPOSX1_1087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_1678_), .Q(csr_gpr_iu_gpr_24__18_) );
	DFFPOSX1 DFFPOSX1_1088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_1679_), .Q(csr_gpr_iu_gpr_24__19_) );
	DFFPOSX1 DFFPOSX1_1089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_1680_), .Q(csr_gpr_iu_gpr_24__20_) );
	DFFPOSX1 DFFPOSX1_1090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_1681_), .Q(csr_gpr_iu_gpr_24__21_) );
	DFFPOSX1 DFFPOSX1_1091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_1682_), .Q(csr_gpr_iu_gpr_24__22_) );
	DFFPOSX1 DFFPOSX1_1092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_1683_), .Q(csr_gpr_iu_gpr_24__23_) );
	DFFPOSX1 DFFPOSX1_1093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_1684_), .Q(csr_gpr_iu_gpr_24__24_) );
	DFFPOSX1 DFFPOSX1_1094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_1685_), .Q(csr_gpr_iu_gpr_24__25_) );
	DFFPOSX1 DFFPOSX1_1095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_1686_), .Q(csr_gpr_iu_gpr_24__26_) );
	DFFPOSX1 DFFPOSX1_1096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_1687_), .Q(csr_gpr_iu_gpr_24__27_) );
	DFFPOSX1 DFFPOSX1_1097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_1688_), .Q(csr_gpr_iu_gpr_24__28_) );
	DFFPOSX1 DFFPOSX1_1098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_1689_), .Q(csr_gpr_iu_gpr_24__29_) );
	DFFPOSX1 DFFPOSX1_1099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_1690_), .Q(csr_gpr_iu_gpr_24__30_) );
	DFFPOSX1 DFFPOSX1_1100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_1691_), .Q(csr_gpr_iu_gpr_24__31_) );
	DFFPOSX1 DFFPOSX1_1101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_1532_), .Q(csr_gpr_iu_gpr_20__0_) );
	DFFPOSX1 DFFPOSX1_1102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_1533_), .Q(csr_gpr_iu_gpr_20__1_) );
	DFFPOSX1 DFFPOSX1_1103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_1534_), .Q(csr_gpr_iu_gpr_20__2_) );
	DFFPOSX1 DFFPOSX1_1104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_1535_), .Q(csr_gpr_iu_gpr_20__3_) );
	DFFPOSX1 DFFPOSX1_1105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_1536_), .Q(csr_gpr_iu_gpr_20__4_) );
	DFFPOSX1 DFFPOSX1_1106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_1537_), .Q(csr_gpr_iu_gpr_20__5_) );
	DFFPOSX1 DFFPOSX1_1107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_1538_), .Q(csr_gpr_iu_gpr_20__6_) );
	DFFPOSX1 DFFPOSX1_1108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_1539_), .Q(csr_gpr_iu_gpr_20__7_) );
	DFFPOSX1 DFFPOSX1_1109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_1540_), .Q(csr_gpr_iu_gpr_20__8_) );
	DFFPOSX1 DFFPOSX1_1110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_1541_), .Q(csr_gpr_iu_gpr_20__9_) );
	DFFPOSX1 DFFPOSX1_1111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_1542_), .Q(csr_gpr_iu_gpr_20__10_) );
	DFFPOSX1 DFFPOSX1_1112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_1543_), .Q(csr_gpr_iu_gpr_20__11_) );
	DFFPOSX1 DFFPOSX1_1113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_1544_), .Q(csr_gpr_iu_gpr_20__12_) );
	DFFPOSX1 DFFPOSX1_1114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_1545_), .Q(csr_gpr_iu_gpr_20__13_) );
	DFFPOSX1 DFFPOSX1_1115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_1546_), .Q(csr_gpr_iu_gpr_20__14_) );
	DFFPOSX1 DFFPOSX1_1116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1547_), .Q(csr_gpr_iu_gpr_20__15_) );
	DFFPOSX1 DFFPOSX1_1117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1548_), .Q(csr_gpr_iu_gpr_20__16_) );
	DFFPOSX1 DFFPOSX1_1118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1549_), .Q(csr_gpr_iu_gpr_20__17_) );
	DFFPOSX1 DFFPOSX1_1119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1550_), .Q(csr_gpr_iu_gpr_20__18_) );
	DFFPOSX1 DFFPOSX1_1120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1551_), .Q(csr_gpr_iu_gpr_20__19_) );
	DFFPOSX1 DFFPOSX1_1121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_1552_), .Q(csr_gpr_iu_gpr_20__20_) );
	DFFPOSX1 DFFPOSX1_1122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1553_), .Q(csr_gpr_iu_gpr_20__21_) );
	DFFPOSX1 DFFPOSX1_1123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1554_), .Q(csr_gpr_iu_gpr_20__22_) );
	DFFPOSX1 DFFPOSX1_1124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1555_), .Q(csr_gpr_iu_gpr_20__23_) );
	DFFPOSX1 DFFPOSX1_1125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1556_), .Q(csr_gpr_iu_gpr_20__24_) );
	DFFPOSX1 DFFPOSX1_1126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1557_), .Q(csr_gpr_iu_gpr_20__25_) );
	DFFPOSX1 DFFPOSX1_1127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1558_), .Q(csr_gpr_iu_gpr_20__26_) );
	DFFPOSX1 DFFPOSX1_1128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_1559_), .Q(csr_gpr_iu_gpr_20__27_) );
	DFFPOSX1 DFFPOSX1_1129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_1560_), .Q(csr_gpr_iu_gpr_20__28_) );
	DFFPOSX1 DFFPOSX1_1130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_1561_), .Q(csr_gpr_iu_gpr_20__29_) );
	DFFPOSX1 DFFPOSX1_1131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_1562_), .Q(csr_gpr_iu_gpr_20__30_) );
	DFFPOSX1 DFFPOSX1_1132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_1563_), .Q(csr_gpr_iu_gpr_20__31_) );
	DFFPOSX1 DFFPOSX1_1133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_2204_), .Q(csr_gpr_iu_gpr_13__0_) );
	DFFPOSX1 DFFPOSX1_1134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_2205_), .Q(csr_gpr_iu_gpr_13__1_) );
	DFFPOSX1 DFFPOSX1_1135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_2206_), .Q(csr_gpr_iu_gpr_13__2_) );
	DFFPOSX1 DFFPOSX1_1136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_2207_), .Q(csr_gpr_iu_gpr_13__3_) );
	DFFPOSX1 DFFPOSX1_1137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_2208_), .Q(csr_gpr_iu_gpr_13__4_) );
	DFFPOSX1 DFFPOSX1_1138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_2209_), .Q(csr_gpr_iu_gpr_13__5_) );
	DFFPOSX1 DFFPOSX1_1139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_2210_), .Q(csr_gpr_iu_gpr_13__6_) );
	DFFPOSX1 DFFPOSX1_1140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_2211_), .Q(csr_gpr_iu_gpr_13__7_) );
	DFFPOSX1 DFFPOSX1_1141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_2212_), .Q(csr_gpr_iu_gpr_13__8_) );
	DFFPOSX1 DFFPOSX1_1142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_2213_), .Q(csr_gpr_iu_gpr_13__9_) );
	DFFPOSX1 DFFPOSX1_1143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_2214_), .Q(csr_gpr_iu_gpr_13__10_) );
	DFFPOSX1 DFFPOSX1_1144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_2215_), .Q(csr_gpr_iu_gpr_13__11_) );
	DFFPOSX1 DFFPOSX1_1145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_2216_), .Q(csr_gpr_iu_gpr_13__12_) );
	DFFPOSX1 DFFPOSX1_1146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_2217_), .Q(csr_gpr_iu_gpr_13__13_) );
	DFFPOSX1 DFFPOSX1_1147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_2218_), .Q(csr_gpr_iu_gpr_13__14_) );
	DFFPOSX1 DFFPOSX1_1148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_2219_), .Q(csr_gpr_iu_gpr_13__15_) );
	DFFPOSX1 DFFPOSX1_1149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_2220_), .Q(csr_gpr_iu_gpr_13__16_) );
	DFFPOSX1 DFFPOSX1_1150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_2221_), .Q(csr_gpr_iu_gpr_13__17_) );
	DFFPOSX1 DFFPOSX1_1151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_2222_), .Q(csr_gpr_iu_gpr_13__18_) );
	DFFPOSX1 DFFPOSX1_1152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_2223_), .Q(csr_gpr_iu_gpr_13__19_) );
	DFFPOSX1 DFFPOSX1_1153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_2224_), .Q(csr_gpr_iu_gpr_13__20_) );
	DFFPOSX1 DFFPOSX1_1154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_2225_), .Q(csr_gpr_iu_gpr_13__21_) );
	DFFPOSX1 DFFPOSX1_1155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_2226_), .Q(csr_gpr_iu_gpr_13__22_) );
	DFFPOSX1 DFFPOSX1_1156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_2227_), .Q(csr_gpr_iu_gpr_13__23_) );
	DFFPOSX1 DFFPOSX1_1157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_2228_), .Q(csr_gpr_iu_gpr_13__24_) );
	DFFPOSX1 DFFPOSX1_1158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_2229_), .Q(csr_gpr_iu_gpr_13__25_) );
	DFFPOSX1 DFFPOSX1_1159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_2230_), .Q(csr_gpr_iu_gpr_13__26_) );
	DFFPOSX1 DFFPOSX1_1160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_2231_), .Q(csr_gpr_iu_gpr_13__27_) );
	DFFPOSX1 DFFPOSX1_1161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_2232_), .Q(csr_gpr_iu_gpr_13__28_) );
	DFFPOSX1 DFFPOSX1_1162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_2233_), .Q(csr_gpr_iu_gpr_13__29_) );
	DFFPOSX1 DFFPOSX1_1163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_2234_), .Q(csr_gpr_iu_gpr_13__30_) );
	DFFPOSX1 DFFPOSX1_1164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_2235_), .Q(csr_gpr_iu_gpr_13__31_) );
	DFFPOSX1 DFFPOSX1_1165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_1467__0_), .Q(biu_exce_chk_statu_cpu_0_) );
	DFFPOSX1 DFFPOSX1_1166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_1467__1_), .Q(biu_exce_chk_statu_cpu_1_) );
	DFFPOSX1 DFFPOSX1_1167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_1467__2_), .Q(biu_exce_chk_statu_cpu_2_) );
	DFFPOSX1 DFFPOSX1_1168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_1467__3_), .Q(biu_exce_chk_statu_cpu_3_) );
	DFFPOSX1 DFFPOSX1_1169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_1459_), .Q(csr_gpr_iu_ins_addr_mis_reg) );
	DFFPOSX1 DFFPOSX1_1170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_1458_), .Q(csr_gpr_iu_ins_acc_fault_reg) );
	DFFPOSX1 DFFPOSX1_1171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_1463_), .Q(csr_gpr_iu_load_addr_mis_reg) );
	DFFPOSX1 DFFPOSX1_1172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_1462_), .Q(csr_gpr_iu_load_acc_fault_reg) );
	DFFPOSX1 DFFPOSX1_1173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_1465_), .Q(csr_gpr_iu_st_addr_mis_reg) );
	DFFPOSX1 DFFPOSX1_1174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_1464_), .Q(csr_gpr_iu_st_acc_fault_reg) );
	DFFPOSX1 DFFPOSX1_1175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_1460_), .Q(csr_gpr_iu_ins_page_fault_reg) );
	DFFPOSX1 DFFPOSX1_1176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_1461_), .Q(csr_gpr_iu_ld_page_fault_reg) );
	DFFPOSX1 DFFPOSX1_1177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_1466_), .Q(csr_gpr_iu_st_page_fault_reg) );
	NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(biu_exce_chk_statu_cpu_0_), .Y(_6756_) );
	NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_2_), .Y(_6757_) );
	INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(_6757_), .Y(_6758_) );
	NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .Y(_6759_) );
	INVX1 INVX1_1126 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_23_), .Y(_6760_) );
	INVX1 INVX1_1127 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_22_), .Y(_6761_) );
	NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_21_), .B(csr_gpr_iu_csr_mcycle_20_), .Y(_6762_) );
	NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_6761_), .C(_6762_), .Y(_6763_) );
	INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_27_), .Y(_6764_) );
	INVX1 INVX1_1128 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_26_), .Y(_6765_) );
	NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_25_), .B(csr_gpr_iu_csr_mcycle_24_), .Y(_6766_) );
	NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6765_), .C(_6766_), .Y(_6767_) );
	NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_6763_), .B(_6767_), .Y(_6768_) );
	NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_29_), .B(csr_gpr_iu_csr_mcycle_28_), .Y(_6769_) );
	NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_31_), .B(csr_gpr_iu_csr_mcycle_30_), .Y(_6770_) );
	AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_6769_), .B(_6770_), .Y(_6771_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_5_), .B(biu_ins_25_bF_buf2), .Y(_6772_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_4_), .B(biu_ins_24_), .Y(_6773_) );
	INVX1 INVX1_1129 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_3_), .Y(_6774_) );
	INVX1 INVX1_1130 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .Y(_6775_) );
	NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_6774_), .B(_6775_), .Y(_6776_) );
	NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_3_), .B(biu_ins_23_), .Y(_6777_) );
	INVX1 INVX1_1131 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_2_), .Y(_6778_) );
	INVX1 INVX1_1132 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf2), .Y(_6779_) );
	NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_6778_), .B(_6779_), .Y(_6780_) );
	NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_2_), .B(biu_ins_22_bF_buf1), .Y(_6781_) );
	AOI22X1 AOI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_6777_), .C(_6780_), .D(_6781_), .Y(_6782_) );
	NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_6772_), .B(_6773_), .C(_6782_), .Y(_6783_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_1_), .B(biu_ins_21_bF_buf0), .Y(_6784_) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_0_), .B(biu_ins_20_bF_buf5), .Y(_6785_) );
	INVX1 INVX1_1133 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_13_), .Y(_6786_) );
	INVX1 INVX1_1134 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_12_), .Y(_6787_) );
	NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_15_), .B(csr_gpr_iu_csr_mcycle_14_), .Y(_6788_) );
	NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_6786_), .B(_6787_), .C(_6788_), .Y(_6789_) );
	INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_19_), .Y(_6790_) );
	INVX1 INVX1_1135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_18_), .Y(_6791_) );
	NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_17_), .B(csr_gpr_iu_csr_mcycle_16_), .Y(_6792_) );
	NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_6790_), .B(_6791_), .C(_6792_), .Y(_6793_) );
	NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_6789_), .B(_6793_), .Y(_6794_) );
	NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .B(_6785_), .C(_6794_), .Y(_6795_) );
	NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_6783_), .B(_6795_), .Y(_6796_) );
	NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_6771_), .C(_6796_), .Y(_6797_) );
	INVX1 INVX1_1136 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_7_), .Y(_6798_) );
	INVX1 INVX1_1137 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf2), .Y(_6799_) );
	NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_6799_), .Y(_6800_) );
	NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_7_), .B(biu_ins_27_bF_buf1), .Y(_6801_) );
	OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(biu_ins_26_bF_buf2), .Y(_6802_) );
	NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(biu_ins_26_bF_buf1), .Y(_6803_) );
	AOI22X1 AOI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_6802_), .B(_6803_), .C(_6800_), .D(_6801_), .Y(_6804_) );
	NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_9_), .B(biu_ins_29_bF_buf2), .Y(_6805_) );
	OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_9_), .B(biu_ins_29_bF_buf1), .Y(_6806_) );
	INVX1 INVX1_1138 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf2), .Y(_6807_) );
	INVX1 INVX1_1139 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_8_), .Y(_6808_) );
	NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_6808_), .Y(_6809_) );
	NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf1), .B(csr_gpr_iu_csr_mcycle_8_), .Y(_6810_) );
	AOI22X1 AOI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_6806_), .B(_6805_), .C(_6809_), .D(_6810_), .Y(_6811_) );
	INVX1 INVX1_1140 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_10_), .Y(_6812_) );
	INVX1 INVX1_1141 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf2), .Y(_6813_) );
	NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_6812_), .B(_6813_), .Y(_6814_) );
	NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_10_), .B(biu_ins_30_bF_buf1), .Y(_6815_) );
	OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_11_), .B(biu_ins_31_bF_buf5), .Y(_6816_) );
	NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_11_), .B(biu_ins_31_bF_buf4), .Y(_6817_) );
	AOI22X1 AOI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_6816_), .B(_6817_), .C(_6814_), .D(_6815_), .Y(_6818_) );
	NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .B(_6811_), .C(_6818_), .Y(_6819_) );
	OAI21X1 OAI21X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .C(_6759__bF_buf4), .Y(_6820_) );
	INVX8 INVX8_54 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf3), .Y(_6821_) );
	INVX1 INVX1_1142 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_0_), .Y(_6822_) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .B(csr_gpr_iu_csr_minstret_4_), .Y(_6823_) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf1), .B(csr_gpr_iu_csr_minstret_5_), .Y(_6824_) );
	OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf0), .B(csr_gpr_iu_csr_minstret_2_), .Y(_6825_) );
	NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf3), .B(csr_gpr_iu_csr_minstret_2_), .Y(_6826_) );
	INVX1 INVX1_1143 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_3_), .Y(_6827_) );
	NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_6775_), .B(_6827_), .Y(_6828_) );
	NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .B(csr_gpr_iu_csr_minstret_3_), .Y(_6829_) );
	AOI22X1 AOI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_6825_), .B(_6826_), .C(_6828_), .D(_6829_), .Y(_6830_) );
	NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_6823_), .B(_6824_), .C(_6830_), .Y(_6831_) );
	INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_15_), .Y(_6832_) );
	INVX1 INVX1_1144 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_14_), .Y(_6833_) );
	NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_13_), .B(csr_gpr_iu_csr_minstret_12_), .Y(_6834_) );
	NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6833_), .C(_6834_), .Y(_6835_) );
	INVX1 INVX1_1145 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_17_), .Y(_6836_) );
	INVX1 INVX1_1146 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_16_), .Y(_6837_) );
	NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_19_), .B(csr_gpr_iu_csr_minstret_18_), .Y(_6838_) );
	NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .B(_6837_), .C(_6838_), .Y(_6839_) );
	NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_6835_), .B(_6839_), .Y(_6840_) );
	XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf4), .B(csr_gpr_iu_csr_minstret_0_), .Y(_6841_) );
	XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf3), .B(csr_gpr_iu_csr_minstret_1_), .Y(_6842_) );
	NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_6842_), .C(_6840_), .Y(_6843_) );
	NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_6831_), .B(_6843_), .Y(_6844_) );
	INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_23_), .Y(_6845_) );
	INVX1 INVX1_1147 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_22_), .Y(_6846_) );
	NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_21_), .B(csr_gpr_iu_csr_minstret_20_), .Y(_6847_) );
	NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6846_), .C(_6847_), .Y(_6848_) );
	INVX1 INVX1_1148 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_27_), .Y(_6849_) );
	INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_26_), .Y(_6850_) );
	NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_25_), .B(csr_gpr_iu_csr_minstret_24_), .Y(_6851_) );
	NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_6850_), .C(_6851_), .Y(_6852_) );
	OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_6848_), .B(_6852_), .Y(_6853_) );
	INVX1 INVX1_1149 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_31_), .Y(_6854_) );
	INVX1 INVX1_1150 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_30_), .Y(_6855_) );
	NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_29_), .B(csr_gpr_iu_csr_minstret_28_), .Y(_6856_) );
	NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_6854_), .B(_6855_), .C(_6856_), .Y(_6857_) );
	NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_6857_), .B(_6853_), .Y(_6858_) );
	AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_6844_), .B(_6858_), .Y(_6859_) );
	NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf0), .B(csr_gpr_iu_csr_minstret_7_), .Y(_6860_) );
	INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_7_), .Y(_6861_) );
	NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_6799_), .B(_6861_), .Y(_6862_) );
	XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf0), .B(csr_gpr_iu_csr_minstret_6_), .Y(_6863_) );
	OAI21X1 OAI21X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_6860_), .B(_6862_), .C(_6863_), .Y(_6864_) );
	XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf0), .B(csr_gpr_iu_csr_minstret_9_), .Y(_6865_) );
	NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf0), .B(csr_gpr_iu_csr_minstret_8_), .Y(_6866_) );
	INVX1 INVX1_1151 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_8_), .Y(_6867_) );
	NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_6867_), .Y(_6868_) );
	OAI21X1 OAI21X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_6868_), .C(_6865_), .Y(_6869_) );
	OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_6864_), .B(_6869_), .Y(_6870_) );
	NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf0), .B(csr_gpr_iu_csr_minstret_10_), .Y(_6871_) );
	INVX1 INVX1_1152 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_10_), .Y(_6872_) );
	NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_6813_), .B(_6872_), .Y(_6873_) );
	XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(csr_gpr_iu_csr_minstret_11_), .Y(_6874_) );
	OAI21X1 OAI21X1_3168 ( .gnd(gnd), .vdd(vdd), .A(_6871_), .B(_6873_), .C(_6874_), .Y(_6875_) );
	NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_6875_), .B(_6870_), .Y(_6876_) );
	NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6859_), .Y(_6877_) );
	MUX2X1 MUX2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_6822_), .B(addr_csr_0_), .S(_6877_), .Y(_6878_) );
	INVX8 INVX8_55 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf65), .Y(_6879_) );
	OAI21X1 OAI21X1_3169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_0_), .B(_6821__bF_buf3), .C(_6879__bF_buf42), .Y(_6880_) );
	AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_6821__bF_buf2), .B(_6878_), .C(_6880_), .Y(_6712__0_) );
	INVX1 INVX1_1153 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_1_), .Y(_6881_) );
	NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_6822_), .B(_6881_), .Y(_6882_) );
	NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_0_), .B(csr_gpr_iu_csr_minstret_1_), .Y(_6883_) );
	OAI21X1 OAI21X1_3170 ( .gnd(gnd), .vdd(vdd), .A(_6882_), .B(_6883_), .C(_6877_), .Y(_6884_) );
	OAI21X1 OAI21X1_3171 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_6877_), .C(_6884_), .Y(_6885_) );
	OAI21X1 OAI21X1_3172 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_1_), .B(_6821__bF_buf1), .C(_6879__bF_buf41), .Y(_6886_) );
	AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_6821__bF_buf0), .B(_6885_), .C(_6886_), .Y(_6712__1_) );
	NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_2_), .B(_6882_), .Y(_6887_) );
	INVX1 INVX1_1154 ( .gnd(gnd), .vdd(vdd), .A(_6887_), .Y(_6888_) );
	NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_2_), .B(_6882_), .Y(_6889_) );
	OAI21X1 OAI21X1_3173 ( .gnd(gnd), .vdd(vdd), .A(_6888_), .B(_6889_), .C(_6877_), .Y(_6890_) );
	OAI21X1 OAI21X1_3174 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_6877_), .C(_6890_), .Y(_6891_) );
	OAI21X1 OAI21X1_3175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_2_), .B(_6821__bF_buf3), .C(_6879__bF_buf40), .Y(_6892_) );
	AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_6821__bF_buf2), .B(_6891_), .C(_6892_), .Y(_6712__2_) );
	INVX8 INVX8_56 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .Y(_6893_) );
	OAI21X1 OAI21X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_6888_), .B(_6893__bF_buf4), .C(_6821__bF_buf1), .Y(_6894_) );
	INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .Y(_6895_) );
	NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6887_), .Y(_6896_) );
	MUX2X1 MUX2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6895_), .S(_6877_), .Y(_6897_) );
	OAI21X1 OAI21X1_3177 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf2), .B(_6897_), .C(_6879__bF_buf39), .Y(_6898_) );
	AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6894_), .C(_6898_), .Y(_6712__3_) );
	INVX1 INVX1_1155 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_4_), .Y(_6899_) );
	OAI21X1 OAI21X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6893__bF_buf3), .C(_6821__bF_buf0), .Y(_6900_) );
	INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .Y(_6901_) );
	NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_4_), .B(_6896_), .Y(_6902_) );
	INVX1 INVX1_1156 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .Y(_6903_) );
	MUX2X1 MUX2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_6903_), .B(_6901_), .S(_6877_), .Y(_6904_) );
	OAI21X1 OAI21X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf1), .B(_6904_), .C(_6879__bF_buf38), .Y(_6905_) );
	AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_6900_), .C(_6905_), .Y(_6712__4_) );
	INVX1 INVX1_1157 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_5_), .Y(_6906_) );
	OAI21X1 OAI21X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_6903_), .B(_6893__bF_buf2), .C(_6821__bF_buf3), .Y(_6907_) );
	INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .Y(_6908_) );
	NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_6906_), .B(_6902_), .Y(_6909_) );
	MUX2X1 MUX2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_6909_), .B(_6908_), .S(_6877_), .Y(_6910_) );
	OAI21X1 OAI21X1_3181 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf0), .B(_6910_), .C(_6879__bF_buf37), .Y(_6911_) );
	AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_6906_), .B(_6907_), .C(_6911_), .Y(_6712__5_) );
	INVX1 INVX1_1158 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_6_), .Y(_6912_) );
	OAI21X1 OAI21X1_3182 ( .gnd(gnd), .vdd(vdd), .A(_6909_), .B(_6893__bF_buf1), .C(_6821__bF_buf2), .Y(_6913_) );
	INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .Y(_6914_) );
	NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_6_), .B(_6909_), .Y(_6915_) );
	INVX1 INVX1_1159 ( .gnd(gnd), .vdd(vdd), .A(_6915_), .Y(_6916_) );
	MUX2X1 MUX2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_6916_), .B(_6914_), .S(_6877_), .Y(_6917_) );
	OAI21X1 OAI21X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf3), .B(_6917_), .C(_6879__bF_buf36), .Y(_6918_) );
	AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .B(_6913_), .C(_6918_), .Y(_6712__6_) );
	OAI21X1 OAI21X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_6916_), .B(_6893__bF_buf0), .C(_6821__bF_buf1), .Y(_6919_) );
	INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .Y(_6920_) );
	NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6915_), .Y(_6921_) );
	MUX2X1 MUX2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_6921_), .B(_6920_), .S(_6877_), .Y(_6922_) );
	OAI21X1 OAI21X1_3185 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf2), .B(_6922_), .C(_6879__bF_buf35), .Y(_6923_) );
	AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6919_), .C(_6923_), .Y(_6712__7_) );
	NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_8_), .B(_6921_), .Y(_6924_) );
	OAI21X1 OAI21X1_3186 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6915_), .C(_6867_), .Y(_6925_) );
	AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_6925_), .Y(_6926_) );
	INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .Y(_6927_) );
	AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf4), .B(_6927_), .C(_6820__bF_buf1), .Y(_6928_) );
	OAI21X1 OAI21X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf3), .B(_6926_), .C(_6928_), .Y(_6929_) );
	INVX8 INVX8_57 ( .gnd(gnd), .vdd(vdd), .A(_6759__bF_buf3), .Y(_6930_) );
	NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .Y(_6931_) );
	OAI21X1 OAI21X1_3188 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf5), .B(_6931__bF_buf3), .C(csr_gpr_iu_csr_minstret_8_), .Y(_6932_) );
	AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_6929_), .B(_6932_), .C(rst_bF_buf64), .Y(_6712__8_) );
	XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(csr_gpr_iu_csr_minstret_9_), .Y(_6933_) );
	INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .Y(_6934_) );
	AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf2), .B(_6934_), .C(_6820__bF_buf0), .Y(_6935_) );
	OAI21X1 OAI21X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf1), .B(_6933_), .C(_6935_), .Y(_6936_) );
	OAI21X1 OAI21X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf4), .B(_6931__bF_buf2), .C(csr_gpr_iu_csr_minstret_9_), .Y(_6937_) );
	AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_6936_), .B(_6937_), .C(rst_bF_buf63), .Y(_6712__9_) );
	INVX1 INVX1_1160 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_9_), .Y(_6938_) );
	NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6924_), .Y(_6939_) );
	NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_10_), .B(_6939_), .Y(_6940_) );
	OAI21X1 OAI21X1_3191 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6924_), .C(_6872_), .Y(_6941_) );
	AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_6940_), .B(_6941_), .Y(_6942_) );
	INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .Y(_6943_) );
	AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf0), .B(_6943_), .C(_6820__bF_buf3), .Y(_6944_) );
	OAI21X1 OAI21X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf4), .B(_6942_), .C(_6944_), .Y(_6945_) );
	OAI21X1 OAI21X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf3), .B(_6931__bF_buf1), .C(csr_gpr_iu_csr_minstret_10_), .Y(_6946_) );
	AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_6945_), .B(_6946_), .C(rst_bF_buf62), .Y(_6712__10_) );
	XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_6940_), .B(csr_gpr_iu_csr_minstret_11_), .Y(_6947_) );
	INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .Y(_6948_) );
	AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf3), .B(_6948_), .C(_6820__bF_buf2), .Y(_6949_) );
	OAI21X1 OAI21X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf2), .B(_6947_), .C(_6949_), .Y(_6950_) );
	OAI21X1 OAI21X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf2), .B(_6931__bF_buf0), .C(csr_gpr_iu_csr_minstret_11_), .Y(_6951_) );
	AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_6950_), .B(_6951_), .C(rst_bF_buf61), .Y(_6712__11_) );
	INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_11_), .Y(_6952_) );
	NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(_6940_), .Y(_6953_) );
	NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_12_), .B(_6953_), .Y(_6954_) );
	INVX1 INVX1_1161 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_12_), .Y(_6955_) );
	OAI21X1 OAI21X1_3196 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(_6940_), .C(_6955_), .Y(_6956_) );
	AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_6956_), .Y(_6957_) );
	INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .Y(_6958_) );
	AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf1), .B(_6958_), .C(_6820__bF_buf1), .Y(_6959_) );
	OAI21X1 OAI21X1_3197 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf0), .B(_6957_), .C(_6959_), .Y(_6960_) );
	OAI21X1 OAI21X1_3198 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf1), .B(_6931__bF_buf3), .C(csr_gpr_iu_csr_minstret_12_), .Y(_6961_) );
	AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_6960_), .B(_6961_), .C(rst_bF_buf60), .Y(_6712__12_) );
	NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .B(_6931__bF_buf2), .Y(_6962_) );
	AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(addr_csr_13_bF_buf1), .C(_6930__bF_buf0), .Y(_6963_) );
	NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf1), .B(_6954_), .Y(_6964_) );
	XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_6964_), .B(csr_gpr_iu_csr_minstret_13_), .Y(_6965_) );
	OAI21X1 OAI21X1_3199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_13_), .B(_6759__bF_buf2), .C(_6879__bF_buf34), .Y(_6966_) );
	AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_6965_), .B(_6963_), .C(_6966_), .Y(_6712__13_) );
	OAI21X1 OAI21X1_3200 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_14_), .B(_6821__bF_buf0), .C(_6879__bF_buf33), .Y(_6967_) );
	INVX1 INVX1_1162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_13_), .Y(_6968_) );
	OAI21X1 OAI21X1_3201 ( .gnd(gnd), .vdd(vdd), .A(_6968_), .B(_6954_), .C(_6833_), .Y(_6969_) );
	NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_6867_), .B(_6938_), .Y(_6970_) );
	NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_6872_), .B(_6952_), .Y(_6971_) );
	AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .B(_6971_), .Y(_6972_) );
	AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_6921_), .B(_6972_), .Y(_6973_) );
	NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_6968_), .B(_6955_), .Y(_6974_) );
	NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_14_), .B(_6974_), .C(_6973_), .Y(_6975_) );
	OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_6975_), .B(_6820__bF_buf0), .Y(_6976_) );
	AOI22X1 AOI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_6893__bF_buf4), .C(_6976_), .D(_6969_), .Y(_6977_) );
	NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_6967_), .B(_6977_), .Y(_6712__14_) );
	INVX1 INVX1_1163 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf1), .Y(_6978_) );
	NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_6978_), .B(_6877_), .Y(_6979_) );
	NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_15_), .B(_6975_), .Y(_6980_) );
	OAI21X1 OAI21X1_3202 ( .gnd(gnd), .vdd(vdd), .A(_6979_), .B(_6980_), .C(_6821__bF_buf3), .Y(_6981_) );
	OAI21X1 OAI21X1_3203 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf3), .B(_6975_), .C(csr_gpr_iu_csr_minstret_15_), .Y(_6982_) );
	AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_6981_), .B(_6982_), .C(rst_bF_buf59), .Y(_6712__15_) );
	NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6976_), .Y(_6983_) );
	NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_16_), .B(_6983_), .Y(_6984_) );
	OAI21X1 OAI21X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6976_), .C(_6837_), .Y(_6985_) );
	NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_6985_), .B(_6984_), .Y(_6986_) );
	NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_6759__bF_buf1), .C(_6962_), .Y(_6987_) );
	AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_6986_), .B(_6987_), .C(rst_bF_buf58), .Y(_6712__16_) );
	INVX1 INVX1_1164 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf1), .Y(_6988_) );
	NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_6930__bF_buf5), .Y(_6989_) );
	AOI22X1 AOI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(_6989_), .C(csr_gpr_iu_csr_minstret_17_), .D(_6984_), .Y(_6990_) );
	OAI21X1 OAI21X1_3205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_17_), .B(_6984_), .C(_6990_), .Y(_6991_) );
	AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_6991_), .B(_6879__bF_buf32), .Y(_6712__17_) );
	NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .B(_6837_), .Y(_6992_) );
	NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_15_), .B(_6992_), .Y(_6993_) );
	NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_6993_), .B(_6975_), .Y(_6994_) );
	NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_18_), .B(_6994_), .Y(_6995_) );
	INVX1 INVX1_1165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_18_), .Y(_6996_) );
	OAI21X1 OAI21X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_6993_), .B(_6975_), .C(_6996_), .Y(_6997_) );
	AOI22X1 AOI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_6893__bF_buf3), .C(_6997_), .D(_6995_), .Y(_6998_) );
	OAI21X1 OAI21X1_3207 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_18_), .B(_6821__bF_buf2), .C(_6879__bF_buf31), .Y(_6999_) );
	AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .B(_6821__bF_buf1), .C(_6999_), .Y(_6712__18_) );
	AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(addr_csr_19_bF_buf1), .C(_6930__bF_buf4), .Y(_7000_) );
	NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf0), .B(_6995_), .Y(_7001_) );
	XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_7001_), .B(csr_gpr_iu_csr_minstret_19_), .Y(_7002_) );
	OAI21X1 OAI21X1_3208 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_19_), .B(_6759__bF_buf0), .C(_6879__bF_buf30), .Y(_7003_) );
	AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_7002_), .B(_7000_), .C(_7003_), .Y(_6712__19_) );
	INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_20_), .Y(_7004_) );
	NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6833_), .Y(_7005_) );
	NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_6974_), .B(_7005_), .C(_6972_), .Y(_7006_) );
	INVX1 INVX1_1166 ( .gnd(gnd), .vdd(vdd), .A(_7006_), .Y(_7007_) );
	AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_6921_), .B(_7007_), .Y(_7008_) );
	AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_19_), .B(csr_gpr_iu_csr_minstret_18_), .Y(_7009_) );
	AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .B(_7009_), .Y(_7010_) );
	NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_7010_), .B(_7008_), .Y(_7011_) );
	XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_7011_), .B(_7004_), .Y(_7012_) );
	AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf2), .B(addr_csr_20_), .C(_6820__bF_buf2), .Y(_7013_) );
	OAI21X1 OAI21X1_3209 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_20_), .B(_6821__bF_buf0), .C(_6879__bF_buf29), .Y(_7014_) );
	AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_7012_), .B(_7013_), .C(_7014_), .Y(_6712__20_) );
	OAI21X1 OAI21X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(csr_gpr_iu_csr_minstret_21_), .Y(_7015_) );
	NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf1), .B(_6893__bF_buf1), .Y(_7016_) );
	NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_7004_), .B(_7011_), .Y(_7017_) );
	XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_7017_), .B(csr_gpr_iu_csr_minstret_21_), .Y(_7018_) );
	AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_7018_), .B(_7016_), .C(_6931__bF_buf3), .Y(_7019_) );
	INVX1 INVX1_1167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_21_), .Y(_7020_) );
	INVX8 INVX8_58 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf2), .Y(_7021_) );
	NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_7020_), .B(_7021__bF_buf4), .Y(_7022_) );
	OAI21X1 OAI21X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7019_), .C(_6759__bF_buf4), .Y(_7023_) );
	AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_7023_), .B(_7015_), .C(rst_bF_buf57), .Y(_6712__21_) );
	NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_7020_), .B(_7004_), .Y(_7024_) );
	INVX1 INVX1_1168 ( .gnd(gnd), .vdd(vdd), .A(_7024_), .Y(_7025_) );
	NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_7011_), .Y(_7026_) );
	XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_7026_), .B(csr_gpr_iu_csr_minstret_22_), .Y(_7027_) );
	AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf0), .B(addr_csr_22_), .C(_6820__bF_buf1), .Y(_7028_) );
	OAI21X1 OAI21X1_3212 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_22_), .B(_6821__bF_buf3), .C(_6879__bF_buf28), .Y(_7029_) );
	AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .B(_7028_), .C(_7029_), .Y(_6712__22_) );
	OAI21X1 OAI21X1_3213 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(csr_gpr_iu_csr_minstret_23_), .Y(_7030_) );
	NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf1), .B(_6893__bF_buf4), .Y(_7031_) );
	AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_7008_), .B(_7010_), .Y(_7032_) );
	NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_22_), .B(_7024_), .C(_7032_), .Y(_7033_) );
	XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_7033_), .B(_6845_), .Y(_7034_) );
	AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_7034_), .B(_7031_), .C(_6931__bF_buf1), .Y(_7035_) );
	NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_7021__bF_buf3), .Y(_7036_) );
	OAI21X1 OAI21X1_3214 ( .gnd(gnd), .vdd(vdd), .A(_7036_), .B(_7035_), .C(_6759__bF_buf3), .Y(_7037_) );
	AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .B(_7030_), .C(rst_bF_buf56), .Y(_6712__23_) );
	INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_24_), .Y(_7038_) );
	NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6846_), .Y(_7039_) );
	NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_7024_), .B(_7039_), .C(_7010_), .Y(_7040_) );
	INVX1 INVX1_1169 ( .gnd(gnd), .vdd(vdd), .A(_7040_), .Y(_7041_) );
	NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_7041_), .B(_7008_), .Y(_7042_) );
	XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_7042_), .B(_7038_), .Y(_7043_) );
	AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf3), .B(addr_csr_24_), .C(_6820__bF_buf0), .Y(_7044_) );
	OAI21X1 OAI21X1_3215 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_24_), .B(_6821__bF_buf2), .C(_6879__bF_buf27), .Y(_7045_) );
	AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_7043_), .B(_7044_), .C(_7045_), .Y(_6712__24_) );
	OAI21X1 OAI21X1_3216 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(csr_gpr_iu_csr_minstret_25_), .Y(_7046_) );
	NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf1), .B(_6893__bF_buf2), .Y(_7047_) );
	NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_7038_), .B(_7042_), .Y(_7048_) );
	XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_7048_), .B(csr_gpr_iu_csr_minstret_25_), .Y(_7049_) );
	AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_7049_), .B(_7047_), .C(_6931__bF_buf0), .Y(_7050_) );
	INVX1 INVX1_1170 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_25_), .Y(_7051_) );
	NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_7051_), .B(_7021__bF_buf2), .Y(_7052_) );
	OAI21X1 OAI21X1_3217 ( .gnd(gnd), .vdd(vdd), .A(_7052_), .B(_7050_), .C(_6759__bF_buf2), .Y(_7053_) );
	AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_7053_), .B(_7046_), .C(rst_bF_buf55), .Y(_6712__25_) );
	NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_7051_), .B(_7038_), .Y(_7054_) );
	NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_7041_), .B(_7054_), .C(_7008_), .Y(_7055_) );
	XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_7055_), .B(_6850_), .Y(_7056_) );
	AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf1), .B(addr_csr_26_), .C(_6820__bF_buf3), .Y(_7057_) );
	OAI21X1 OAI21X1_3218 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_26_), .B(_6821__bF_buf1), .C(_6879__bF_buf26), .Y(_7058_) );
	AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_7056_), .B(_7057_), .C(_7058_), .Y(_6712__26_) );
	OAI21X1 OAI21X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(csr_gpr_iu_csr_minstret_27_), .Y(_7059_) );
	NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf1), .B(_6893__bF_buf0), .Y(_7060_) );
	OAI21X1 OAI21X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_7055_), .C(csr_gpr_iu_csr_minstret_27_), .Y(_7061_) );
	NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_7055_), .Y(_7062_) );
	NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_7062_), .Y(_7063_) );
	NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .B(_7061_), .C(_7063_), .Y(_7064_) );
	MUX2X1 MUX2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_7064_), .B(csr_gpr_iu_csr_minstret_27_), .S(_7021__bF_buf1), .Y(_7065_) );
	OAI21X1 OAI21X1_3221 ( .gnd(gnd), .vdd(vdd), .A(_6930__bF_buf3), .B(_7065_), .C(_7059_), .Y(_7066_) );
	AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_6879__bF_buf25), .Y(_6712__27_) );
	INVX1 INVX1_1171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_28_), .Y(_7067_) );
	NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_6850_), .Y(_7068_) );
	AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_7054_), .B(_7068_), .Y(_7069_) );
	INVX1 INVX1_1172 ( .gnd(gnd), .vdd(vdd), .A(_7069_), .Y(_7070_) );
	NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .B(_7070_), .C(_7042_), .Y(_7071_) );
	INVX1 INVX1_1173 ( .gnd(gnd), .vdd(vdd), .A(_7071_), .Y(_7072_) );
	OAI21X1 OAI21X1_3222 ( .gnd(gnd), .vdd(vdd), .A(_7070_), .B(_7042_), .C(_7067_), .Y(_7073_) );
	NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .B(_7072_), .Y(_7074_) );
	AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf4), .B(addr_csr_28_), .C(_6820__bF_buf2), .Y(_7075_) );
	OAI21X1 OAI21X1_3223 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_28_), .B(_6821__bF_buf0), .C(_6879__bF_buf24), .Y(_7076_) );
	AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_7074_), .B(_7075_), .C(_7076_), .Y(_6712__28_) );
	AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(addr_csr_29_bF_buf1), .C(_6930__bF_buf2), .Y(_7077_) );
	OAI21X1 OAI21X1_3224 ( .gnd(gnd), .vdd(vdd), .A(_6797_), .B(_6819_), .C(_7071_), .Y(_7078_) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_7078_), .B(csr_gpr_iu_csr_minstret_29_), .Y(_7079_) );
	OAI21X1 OAI21X1_3225 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_29_), .B(_6759__bF_buf1), .C(_6879__bF_buf23), .Y(_7080_) );
	AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_7079_), .B(_7077_), .C(_7080_), .Y(_6712__29_) );
	NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_29_), .B(_7071_), .Y(_7081_) );
	OAI21X1 OAI21X1_3226 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf1), .B(_7081_), .C(csr_gpr_iu_csr_minstret_30_), .Y(_7082_) );
	NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_6820__bF_buf0), .B(_7081_), .Y(_7083_) );
	INVX1 INVX1_1174 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .Y(_7084_) );
	NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_6930__bF_buf1), .Y(_7085_) );
	AOI22X1 AOI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(_7085_), .C(_6855_), .D(_7083_), .Y(_7086_) );
	AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_7086_), .B(_7082_), .C(rst_bF_buf54), .Y(_6712__30_) );
	AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_6893__bF_buf3), .B(addr_csr_31_bF_buf1), .C(_6820__bF_buf3), .Y(_7087_) );
	NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_7081_), .Y(_7088_) );
	XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_7088_), .B(csr_gpr_iu_csr_minstret_31_), .Y(_7089_) );
	OAI21X1 OAI21X1_3227 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_31_), .B(_6821__bF_buf3), .C(_6879__bF_buf22), .Y(_7090_) );
	AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_7089_), .B(_7087_), .C(_7090_), .Y(_6712__31_) );
	INVX1 INVX1_1175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_0_), .Y(_7091_) );
	OAI21X1 OAI21X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(_7091_), .Y(_7092_) );
	OAI21X1 OAI21X1_3229 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_7021__bF_buf0), .C(_6759__bF_buf0), .Y(_7093_) );
	OAI21X1 OAI21X1_3230 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_0_), .B(_6820__bF_buf2), .C(_6879__bF_buf21), .Y(_7094_) );
	AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_7093_), .B(_7092_), .C(_7094_), .Y(_6705__0_) );
	INVX1 INVX1_1176 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_1_), .Y(_7095_) );
	OAI21X1 OAI21X1_3231 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .C(_7095_), .Y(_7096_) );
	OAI21X1 OAI21X1_3232 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_7021__bF_buf4), .C(_7096_), .Y(_7097_) );
	NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_7091_), .B(_7095_), .Y(_7098_) );
	NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_0_), .B(csr_gpr_iu_csr_mcycle_1_), .Y(_7099_) );
	NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_7099_), .B(_7098_), .Y(_7100_) );
	OAI21X1 OAI21X1_3233 ( .gnd(gnd), .vdd(vdd), .A(_6759__bF_buf4), .B(_7100_), .C(_6879__bF_buf20), .Y(_7101_) );
	AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_7097_), .B(_6759__bF_buf3), .C(_7101_), .Y(_6705__1_) );
	OAI21X1 OAI21X1_3234 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .C(_6778_), .Y(_7102_) );
	OAI21X1 OAI21X1_3235 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_7021__bF_buf3), .C(_7102_), .Y(_7103_) );
	NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_2_), .B(_7098_), .Y(_7104_) );
	INVX1 INVX1_1177 ( .gnd(gnd), .vdd(vdd), .A(_7104_), .Y(_7105_) );
	OAI21X1 OAI21X1_3236 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_2_), .B(_7098_), .C(_6930__bF_buf0), .Y(_7106_) );
	OAI22X1 OAI22X1_645 ( .gnd(gnd), .vdd(vdd), .A(_7105_), .B(_7106_), .C(_6930__bF_buf5), .D(_7103_), .Y(_7107_) );
	AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_7107_), .B(_6879__bF_buf19), .Y(_6705__2_) );
	NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_6774_), .B(_7104_), .Y(_7108_) );
	OAI21X1 OAI21X1_3237 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_3_), .B(_7105_), .C(_6930__bF_buf4), .Y(_7109_) );
	AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_7021__bF_buf2), .B(_6774_), .C(_6930__bF_buf3), .Y(_7110_) );
	OAI21X1 OAI21X1_3238 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_7021__bF_buf1), .C(_7110_), .Y(_7111_) );
	OAI21X1 OAI21X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .B(_7109_), .C(_7111_), .Y(_7112_) );
	AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_7112_), .B(_6879__bF_buf18), .Y(_6705__3_) );
	NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_4_), .B(_7108_), .Y(_7113_) );
	INVX1 INVX1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7113_), .Y(_7114_) );
	OAI21X1 OAI21X1_3240 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_4_), .B(_7108_), .C(_6930__bF_buf2), .Y(_7115_) );
	OAI21X1 OAI21X1_3241 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .C(csr_gpr_iu_csr_mcycle_4_), .Y(_7116_) );
	OAI21X1 OAI21X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_7021__bF_buf0), .C(_7116_), .Y(_7117_) );
	NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_6759__bF_buf2), .B(_7117_), .Y(_7118_) );
	OAI21X1 OAI21X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_7114_), .B(_7115_), .C(_7118_), .Y(_7119_) );
	AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_7119_), .B(_6879__bF_buf17), .Y(_6705__4_) );
	INVX1 INVX1_1179 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_5_), .Y(_7120_) );
	OAI21X1 OAI21X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6797_), .C(_7120_), .Y(_7121_) );
	OAI21X1 OAI21X1_3245 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_7021__bF_buf4), .C(_7121_), .Y(_7122_) );
	NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_5_), .B(_7114_), .Y(_7123_) );
	NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_7120_), .B(_7113_), .Y(_7124_) );
	OAI21X1 OAI21X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(_7123_), .C(_6930__bF_buf1), .Y(_7125_) );
	NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf16), .B(_7125_), .Y(_7126_) );
	AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .B(_6759__bF_buf1), .C(_7126_), .Y(_6705__5_) );
	NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(_7124_), .Y(_7127_) );
	INVX1 INVX1_1180 ( .gnd(gnd), .vdd(vdd), .A(_7127_), .Y(_7128_) );
	OAI21X1 OAI21X1_3247 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(_7124_), .C(_6930__bF_buf0), .Y(_7129_) );
	NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_7021__bF_buf3), .Y(_7130_) );
	OAI21X1 OAI21X1_3248 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(_6931__bF_buf3), .C(_6759__bF_buf0), .Y(_7131_) );
	OAI22X1 OAI22X1_646 ( .gnd(gnd), .vdd(vdd), .A(_7128_), .B(_7129_), .C(_7131_), .D(_7130_), .Y(_7132_) );
	AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_7132_), .B(_6879__bF_buf15), .Y(_6705__6_) );
	NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_7127_), .Y(_7133_) );
	OAI21X1 OAI21X1_3249 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_7_), .B(_7128_), .C(_6930__bF_buf5), .Y(_7134_) );
	AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_7021__bF_buf2), .B(_6798_), .C(_6930__bF_buf4), .Y(_7135_) );
	OAI21X1 OAI21X1_3250 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_7021__bF_buf1), .C(_7135_), .Y(_7136_) );
	OAI21X1 OAI21X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7134_), .C(_7136_), .Y(_7137_) );
	AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_7137_), .B(_6879__bF_buf14), .Y(_6705__7_) );
	NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_8_), .B(_7133_), .Y(_7138_) );
	INVX1 INVX1_1181 ( .gnd(gnd), .vdd(vdd), .A(_7138_), .Y(_7139_) );
	OAI21X1 OAI21X1_3252 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_8_), .B(_7133_), .C(_6930__bF_buf3), .Y(_7140_) );
	AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_7021__bF_buf0), .B(_6808_), .C(_6930__bF_buf2), .Y(_7141_) );
	OAI21X1 OAI21X1_3253 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_7021__bF_buf4), .C(_7141_), .Y(_7142_) );
	OAI21X1 OAI21X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_7139_), .B(_7140_), .C(_7142_), .Y(_7143_) );
	AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_7143_), .B(_6879__bF_buf13), .Y(_6705__8_) );
	AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf2), .B(_6934_), .C(_6930__bF_buf1), .Y(_7144_) );
	OAI21X1 OAI21X1_3255 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_9_), .B(_6931__bF_buf1), .C(_7144_), .Y(_7145_) );
	INVX1 INVX1_1182 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .Y(_7146_) );
	NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_8_), .B(csr_gpr_iu_csr_mcycle_9_), .Y(_7147_) );
	NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7146_), .Y(_7148_) );
	NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_6759__bF_buf4), .B(_7148_), .Y(_7149_) );
	OAI21X1 OAI21X1_3256 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_9_), .B(_7139_), .C(_7149_), .Y(_7150_) );
	AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_7150_), .B(_7145_), .C(rst_bF_buf53), .Y(_6705__9_) );
	NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_10_), .B(_7148_), .Y(_7151_) );
	INVX1 INVX1_1183 ( .gnd(gnd), .vdd(vdd), .A(_7151_), .Y(_7152_) );
	OAI21X1 OAI21X1_3257 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_10_), .B(_7148_), .C(_6930__bF_buf0), .Y(_7153_) );
	AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_7021__bF_buf3), .B(_6812_), .C(_6930__bF_buf5), .Y(_7154_) );
	OAI21X1 OAI21X1_3258 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_7021__bF_buf2), .C(_7154_), .Y(_7155_) );
	OAI21X1 OAI21X1_3259 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .B(_7152_), .C(_7155_), .Y(_7156_) );
	AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_7156_), .B(_6879__bF_buf12), .Y(_6705__10_) );
	AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf0), .B(_6948_), .C(_6930__bF_buf4), .Y(_7157_) );
	OAI21X1 OAI21X1_3260 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_11_), .B(_6931__bF_buf3), .C(_7157_), .Y(_7158_) );
	NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_10_), .B(csr_gpr_iu_csr_mcycle_11_), .Y(_7159_) );
	NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7159_), .Y(_7160_) );
	NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .B(_7133_), .Y(_7161_) );
	OAI21X1 OAI21X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(_7161_), .Y(_7162_) );
	INVX1 INVX1_1184 ( .gnd(gnd), .vdd(vdd), .A(_7162_), .Y(_7163_) );
	OAI21X1 OAI21X1_3262 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_11_), .B(_7152_), .C(_7163_), .Y(_7164_) );
	AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_7164_), .B(_7158_), .C(rst_bF_buf52), .Y(_6705__11_) );
	OAI21X1 OAI21X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_7021__bF_buf1), .C(_6759__bF_buf3), .Y(_7165_) );
	NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_7162_), .B(_7165_), .Y(_7166_) );
	NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(_7161_), .Y(_7167_) );
	OAI21X1 OAI21X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6758_), .C(_7167_), .Y(_7168_) );
	NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf11), .B(_7168_), .Y(_7169_) );
	AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(_7166_), .C(_7169_), .Y(_6705__12_) );
	NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_6786_), .B(_7168_), .Y(_7170_) );
	INVX1 INVX1_1185 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .Y(_7171_) );
	NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf0), .B(_6759__bF_buf2), .Y(_7172_) );
	OAI21X1 OAI21X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_7172_), .B(_7021__bF_buf0), .C(_6786_), .Y(_7173_) );
	OAI21X1 OAI21X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_7173_), .B(_7171_), .C(_6879__bF_buf10), .Y(_7174_) );
	NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_7170_), .B(_7174_), .Y(_6705__13_) );
	INVX1 INVX1_1186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_14_), .Y(_7175_) );
	NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_6759__bF_buf1), .Y(_7176_) );
	OAI21X1 OAI21X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_7176_), .B(_7021__bF_buf4), .C(_7175_), .Y(_7177_) );
	OAI21X1 OAI21X1_3268 ( .gnd(gnd), .vdd(vdd), .A(_7177_), .B(_7170_), .C(_6879__bF_buf9), .Y(_7178_) );
	AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_14_), .B(_7170_), .C(_7178_), .Y(_6705__14_) );
	NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_14_), .B(_7170_), .Y(_7179_) );
	NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_6978_), .B(_6930__bF_buf3), .Y(_7180_) );
	AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf2), .B(_7180_), .C(csr_gpr_iu_csr_mcycle_15_), .Y(_7181_) );
	NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_13_), .B(csr_gpr_iu_csr_mcycle_15_), .C(csr_gpr_iu_csr_mcycle_14_), .Y(_7182_) );
	OAI21X1 OAI21X1_3269 ( .gnd(gnd), .vdd(vdd), .A(_7182_), .B(_7168_), .C(_6879__bF_buf8), .Y(_7183_) );
	AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .B(_7181_), .C(_7183_), .Y(_6705__15_) );
	NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_7182_), .B(_7168_), .Y(_7184_) );
	INVX1 INVX1_1187 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_16_), .Y(_7185_) );
	NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_6759__bF_buf0), .Y(_7186_) );
	OAI21X1 OAI21X1_3270 ( .gnd(gnd), .vdd(vdd), .A(_7186_), .B(_7021__bF_buf3), .C(_7185_), .Y(_7187_) );
	OAI21X1 OAI21X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_7187_), .B(_7184_), .C(_6879__bF_buf7), .Y(_7188_) );
	AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_16_), .B(_7184_), .C(_7188_), .Y(_6705__16_) );
	NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_16_), .B(_7184_), .Y(_7189_) );
	AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf1), .B(_6989_), .C(csr_gpr_iu_csr_mcycle_17_), .Y(_7190_) );
	INVX1 INVX1_1188 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_17_), .Y(_7191_) );
	NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_7191_), .B(_7185_), .Y(_7192_) );
	NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7184_), .Y(_7193_) );
	NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf6), .B(_7193_), .Y(_7194_) );
	AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_7189_), .B(_7190_), .C(_7194_), .Y(_6705__17_) );
	INVX1 INVX1_1189 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .Y(_7195_) );
	NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_7182_), .B(_7195_), .Y(_7196_) );
	INVX1 INVX1_1190 ( .gnd(gnd), .vdd(vdd), .A(_7196_), .Y(_7197_) );
	NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_7197_), .B(_7168_), .Y(_7198_) );
	NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_6759__bF_buf4), .Y(_7199_) );
	OAI21X1 OAI21X1_3272 ( .gnd(gnd), .vdd(vdd), .A(_7199_), .B(_7021__bF_buf2), .C(_6791_), .Y(_7200_) );
	OAI21X1 OAI21X1_3273 ( .gnd(gnd), .vdd(vdd), .A(_7200_), .B(_7198_), .C(_6879__bF_buf5), .Y(_7201_) );
	NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_6791_), .B(_7193_), .Y(_7202_) );
	NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_7201_), .B(_7202_), .Y(_6705__18_) );
	NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_6790_), .B(_6791_), .Y(_7203_) );
	NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_7203_), .B(_7196_), .Y(_7204_) );
	NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .B(_7168_), .Y(_7205_) );
	NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf0), .B(_6759__bF_buf3), .Y(_7206_) );
	OAI21X1 OAI21X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_7206_), .B(_7021__bF_buf1), .C(_6790_), .Y(_7207_) );
	OAI21X1 OAI21X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_7207_), .B(_7202_), .C(_6879__bF_buf4), .Y(_7208_) );
	NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_7205_), .B(_7208_), .Y(_6705__19_) );
	NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_20_), .B(_7203_), .Y(_7209_) );
	INVX1 INVX1_1191 ( .gnd(gnd), .vdd(vdd), .A(_7209_), .Y(_7210_) );
	AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_7198_), .B(_7210_), .Y(_7211_) );
	INVX1 INVX1_1192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_20_), .Y(_7212_) );
	NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_6759__bF_buf2), .Y(_7213_) );
	OAI21X1 OAI21X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .B(_7021__bF_buf0), .C(_7212_), .Y(_7214_) );
	OAI21X1 OAI21X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(_7205_), .C(_6879__bF_buf3), .Y(_7215_) );
	NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_7211_), .B(_7215_), .Y(_6705__20_) );
	INVX1 INVX1_1193 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_21_), .Y(_7216_) );
	NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf0), .B(_6759__bF_buf1), .Y(_7217_) );
	OAI21X1 OAI21X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_7217_), .B(_7021__bF_buf4), .C(_7216_), .Y(_7218_) );
	OAI21X1 OAI21X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_7218_), .B(_7211_), .C(_6879__bF_buf2), .Y(_7219_) );
	AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_21_), .B(_7211_), .C(_7219_), .Y(_6705__21_) );
	NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_7216_), .B(_7212_), .Y(_7220_) );
	NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_6759__bF_buf0), .Y(_7221_) );
	OAI21X1 OAI21X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_7221_), .B(_7021__bF_buf3), .C(_6761_), .Y(_7222_) );
	AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_7205_), .B(_7220_), .C(_7222_), .Y(_7223_) );
	NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_22_), .B(_7220_), .C(_7205_), .Y(_7224_) );
	NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf1), .B(_7224_), .Y(_7225_) );
	NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_7223_), .B(_7225_), .Y(_6705__22_) );
	INVX1 INVX1_1194 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf0), .Y(_7226_) );
	NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_6930__bF_buf2), .Y(_7227_) );
	AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf0), .B(_7227_), .C(csr_gpr_iu_csr_mcycle_23_), .Y(_7228_) );
	OAI21X1 OAI21X1_3281 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_7224_), .C(_6879__bF_buf0), .Y(_7229_) );
	AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_7224_), .B(_7228_), .C(_7229_), .Y(_6705__23_) );
	NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_22_), .B(_7220_), .Y(_7230_) );
	NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_7230_), .Y(_7231_) );
	INVX1 INVX1_1195 ( .gnd(gnd), .vdd(vdd), .A(_7231_), .Y(_7232_) );
	NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .B(_7232_), .Y(_7233_) );
	AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_7171_), .B(_7233_), .Y(_7234_) );
	AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_7234_), .B(csr_gpr_iu_csr_mcycle_24_), .Y(_7235_) );
	INVX1 INVX1_1196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_24_), .Y(_7236_) );
	NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_6759__bF_buf4), .Y(_7237_) );
	OAI21X1 OAI21X1_3282 ( .gnd(gnd), .vdd(vdd), .A(_7237_), .B(_7021__bF_buf2), .C(_7236_), .Y(_7238_) );
	OAI21X1 OAI21X1_3283 ( .gnd(gnd), .vdd(vdd), .A(_7238_), .B(_7234_), .C(_6879__bF_buf42), .Y(_7239_) );
	NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_7235_), .B(_7239_), .Y(_6705__24_) );
	INVX1 INVX1_1197 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_25_), .Y(_7240_) );
	NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf0), .B(_6759__bF_buf3), .Y(_7241_) );
	OAI21X1 OAI21X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_7241_), .B(_7021__bF_buf1), .C(_7240_), .Y(_7242_) );
	OAI21X1 OAI21X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_7242_), .B(_7235_), .C(_6879__bF_buf41), .Y(_7243_) );
	AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_25_), .B(_7235_), .C(_7243_), .Y(_6705__25_) );
	NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_25_), .B(csr_gpr_iu_csr_mcycle_24_), .C(_7233_), .Y(_7244_) );
	NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_7244_), .B(_7168_), .Y(_7245_) );
	NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .B(_6759__bF_buf2), .Y(_7246_) );
	OAI21X1 OAI21X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_7246_), .B(_7021__bF_buf0), .C(_6765_), .Y(_7247_) );
	OAI21X1 OAI21X1_3287 ( .gnd(gnd), .vdd(vdd), .A(_7247_), .B(_7245_), .C(_6879__bF_buf40), .Y(_7248_) );
	AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_26_), .B(_7245_), .C(_7248_), .Y(_6705__26_) );
	NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_26_), .B(_7245_), .Y(_7249_) );
	NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf0), .B(_6759__bF_buf1), .C(_6931__bF_buf3), .Y(_7250_) );
	AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_7250_), .B(_6764_), .Y(_7251_) );
	AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_7249_), .B(_7251_), .C(rst_bF_buf51), .Y(_7252_) );
	OAI21X1 OAI21X1_3288 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_7249_), .C(_7252_), .Y(_7253_) );
	INVX1 INVX1_1198 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .Y(_6705__27_) );
	NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6765_), .Y(_7254_) );
	INVX1 INVX1_1199 ( .gnd(gnd), .vdd(vdd), .A(_7254_), .Y(_7255_) );
	NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_7255_), .B(_7244_), .Y(_7256_) );
	INVX1 INVX1_1200 ( .gnd(gnd), .vdd(vdd), .A(_7256_), .Y(_7257_) );
	NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_7257_), .B(_7168_), .Y(_7258_) );
	INVX1 INVX1_1201 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_28_), .Y(_7259_) );
	NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_6759__bF_buf0), .Y(_7260_) );
	OAI21X1 OAI21X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(_7021__bF_buf4), .C(_7259_), .Y(_7261_) );
	OAI21X1 OAI21X1_3290 ( .gnd(gnd), .vdd(vdd), .A(_7261_), .B(_7258_), .C(_6879__bF_buf39), .Y(_7262_) );
	AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_28_), .B(_7258_), .C(_7262_), .Y(_6705__28_) );
	INVX1 INVX1_1202 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_29_), .Y(_7263_) );
	NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_28_), .B(_7258_), .Y(_7264_) );
	NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf0), .B(_6759__bF_buf4), .C(_6931__bF_buf2), .Y(_7265_) );
	AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_7265_), .B(_7263_), .Y(_7266_) );
	AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_7264_), .B(_7266_), .C(rst_bF_buf50), .Y(_7267_) );
	OAI21X1 OAI21X1_3291 ( .gnd(gnd), .vdd(vdd), .A(_7263_), .B(_7264_), .C(_7267_), .Y(_7268_) );
	INVX1 INVX1_1203 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .Y(_6705__29_) );
	INVX1 INVX1_1204 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_30_), .Y(_7269_) );
	NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_29_), .B(csr_gpr_iu_csr_mcycle_28_), .C(_6930__bF_buf1), .Y(_7270_) );
	NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_7270_), .B(_7257_), .Y(_7271_) );
	NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .B(_7271_), .Y(_7272_) );
	NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .B(_7272_), .Y(_7273_) );
	INVX1 INVX1_1205 ( .gnd(gnd), .vdd(vdd), .A(_7272_), .Y(_7274_) );
	INVX1 INVX1_1206 ( .gnd(gnd), .vdd(vdd), .A(_7085_), .Y(_7275_) );
	OAI21X1 OAI21X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_7275_), .B(_7021__bF_buf3), .C(_7269_), .Y(_7276_) );
	OAI21X1 OAI21X1_3293 ( .gnd(gnd), .vdd(vdd), .A(_7276_), .B(_7274_), .C(_6879__bF_buf38), .Y(_7277_) );
	NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_7273_), .B(_7277_), .Y(_6705__30_) );
	INVX1 INVX1_1207 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf0), .Y(_7278_) );
	NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_7278_), .B(_6930__bF_buf0), .Y(_7279_) );
	AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_6931__bF_buf1), .B(_7279_), .C(csr_gpr_iu_csr_mcycle_31_), .Y(_7280_) );
	OAI21X1 OAI21X1_3294 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .B(_7272_), .C(_7280_), .Y(_7281_) );
	NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_31_), .B(_7273_), .Y(_7282_) );
	NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf37), .B(_7281_), .C(_7282_), .Y(_7283_) );
	INVX1 INVX1_1208 ( .gnd(gnd), .vdd(vdd), .A(_7283_), .Y(_6705__31_) );
	INVX1 INVX1_1209 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_ssip), .Y(_7284_) );
	INVX1 INVX1_1210 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7285_) );
	OAI21X1 OAI21X1_3295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_ssip_in), .B(_7285_), .C(_6879__bF_buf36), .Y(_7286_) );
	AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_7284_), .B(_7285_), .C(_7286_), .Y(_6748_) );
	INVX1 INVX1_1211 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_msip), .Y(_7287_) );
	INVX1 INVX1_1212 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7288_) );
	OAI21X1 OAI21X1_3296 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_msip_in), .B(_7288_), .C(_6879__bF_buf35), .Y(_7289_) );
	AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_7287_), .B(_7288_), .C(_7289_), .Y(_6718_) );
	INVX1 INVX1_1213 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stip), .Y(_7290_) );
	INVX1 INVX1_1214 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7291_) );
	OAI21X1 OAI21X1_3297 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stip_in), .B(_7291_), .C(_6879__bF_buf34), .Y(_7292_) );
	AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_7291_), .C(_7292_), .Y(_6750_) );
	INVX1 INVX1_1215 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtip), .Y(_7293_) );
	INVX1 INVX1_1216 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7294_) );
	OAI21X1 OAI21X1_3298 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtip_in), .B(_7294_), .C(_6879__bF_buf33), .Y(_7295_) );
	AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_7293_), .B(_7294_), .C(_7295_), .Y(_6721_) );
	INVX1 INVX1_1217 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seip), .Y(_7296_) );
	INVX1 INVX1_1218 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7297_) );
	OAI21X1 OAI21X1_3299 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seip_in), .B(_7297_), .C(_6879__bF_buf32), .Y(_7298_) );
	AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_7296_), .B(_7297_), .C(_7298_), .Y(_6741_) );
	INVX1 INVX1_1219 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip), .Y(_7299_) );
	INVX1 INVX1_1220 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_wr), .Y(_7300_) );
	OAI21X1 OAI21X1_3300 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_in), .B(_7300_), .C(_6879__bF_buf31), .Y(_7301_) );
	AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_7299_), .B(_7300_), .C(_7301_), .Y(_6708_) );
	INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_csr_wr), .Y(_7302_) );
	NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf5), .Y(_7303_) );
	INVX8 INVX8_59 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14_bF_buf3), .Y(_7304_) );
	OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf3), .B(biu_ins_31_bF_buf2), .Y(_7305_) );
	NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_7305_), .Y(_7306_) );
	INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(_7306_), .Y(_7307_) );
	NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf3), .B(_7307_), .Y(_7308_) );
	INVX8 INVX8_60 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .Y(_7309_) );
	NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf2), .B(biu_ins_23_), .Y(_7310_) );
	NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf3), .B(biu_ins_21_bF_buf2), .Y(_7311_) );
	NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_7310_), .B(_7311_), .Y(_7312_) );
	INVX1 INVX1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .Y(_7313_) );
	NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .B(biu_ins_25_bF_buf0), .Y(_7314_) );
	INVX1 INVX1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .Y(_7315_) );
	NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf3), .B(_6799_), .Y(_7316_) );
	NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_7316_), .B(_7315_), .Y(_7317_) );
	NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_7313_), .B(_7317_), .Y(_7318_) );
	NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_7318_), .B(_7309__bF_buf3), .Y(_7319_) );
	INVX8 INVX8_61 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .Y(_7320_) );
	OAI21X1 OAI21X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf3), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_0_), .Y(_7321_) );
	NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7308_), .Y(_7322_) );
	NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7322_), .Y(_7323_) );
	INVX1 INVX1_1223 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .Y(_7324_) );
	NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_7324_), .B(_7304__bF_buf13_bF_buf3), .Y(_7325_) );
	NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf3), .B(_7325_), .Y(_7326_) );
	AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_7321_), .B(_7326_), .C(rst_bF_buf49), .Y(_6746__0_) );
	OAI21X1 OAI21X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf3), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_1_), .Y(_7327_) );
	INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .Y(_7328_) );
	NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_7304__bF_buf11_bF_buf3), .Y(_7329_) );
	NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf2), .B(_7329_), .Y(_7330_) );
	AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_7327_), .B(_7330_), .C(rst_bF_buf48), .Y(_6746__1_) );
	OAI21X1 OAI21X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf3), .B(_7320__bF_buf1), .C(csr_gpr_iu_csr_sscratch_2_), .Y(_7331_) );
	INVX1 INVX1_1224 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .Y(_7332_) );
	NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7304__bF_buf9_bF_buf3), .Y(_7333_) );
	NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf1), .B(_7333_), .Y(_7334_) );
	AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_7331_), .B(_7334_), .C(rst_bF_buf47), .Y(_6746__2_) );
	OAI21X1 OAI21X1_3304 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf3), .B(_7320__bF_buf0), .C(csr_gpr_iu_csr_sscratch_3_), .Y(_7335_) );
	NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_6895_), .B(_7304__bF_buf7_bF_buf3), .Y(_7336_) );
	NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf0), .B(_7336_), .Y(_7337_) );
	AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_7335_), .B(_7337_), .C(rst_bF_buf46), .Y(_6746__3_) );
	OAI21X1 OAI21X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf3), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_4_), .Y(_7338_) );
	NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_7304__bF_buf5), .Y(_7339_) );
	NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf3), .B(_7339_), .Y(_7340_) );
	AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_7338_), .B(_7340_), .C(rst_bF_buf45), .Y(_6746__4_) );
	OAI21X1 OAI21X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_5_), .Y(_7341_) );
	NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_7304__bF_buf3), .Y(_7342_) );
	NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf2), .B(_7342_), .Y(_7343_) );
	AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_7341_), .B(_7343_), .C(rst_bF_buf44), .Y(_6746__5_) );
	OAI21X1 OAI21X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_7320__bF_buf1), .C(csr_gpr_iu_csr_sscratch_6_), .Y(_7344_) );
	NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_7304__bF_buf1), .Y(_7345_) );
	NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf1), .B(_7345_), .Y(_7346_) );
	AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_7344_), .B(_7346_), .C(rst_bF_buf43), .Y(_6746__6_) );
	OAI21X1 OAI21X1_3308 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(_7320__bF_buf0), .C(csr_gpr_iu_csr_sscratch_7_), .Y(_7347_) );
	NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_7304__bF_buf14_bF_buf2), .Y(_7348_) );
	NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf0), .B(_7348_), .Y(_7349_) );
	AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_7347_), .B(_7349_), .C(rst_bF_buf42), .Y(_6746__7_) );
	OAI21X1 OAI21X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf2), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_8_), .Y(_7350_) );
	NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_6927_), .B(_7304__bF_buf12_bF_buf2), .Y(_7351_) );
	NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf3), .B(_7351_), .Y(_7352_) );
	AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_7350_), .B(_7352_), .C(rst_bF_buf41), .Y(_6746__8_) );
	OAI21X1 OAI21X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf2), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_9_), .Y(_7353_) );
	NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_7304__bF_buf10_bF_buf2), .Y(_7354_) );
	NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf2), .B(_7354_), .Y(_7355_) );
	AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_7353_), .B(_7355_), .C(rst_bF_buf40), .Y(_6746__9_) );
	OAI21X1 OAI21X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf2), .B(_7320__bF_buf1), .C(csr_gpr_iu_csr_sscratch_10_), .Y(_7356_) );
	NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_7304__bF_buf8_bF_buf2), .Y(_7357_) );
	NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf1), .B(_7357_), .Y(_7358_) );
	AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_7356_), .B(_7358_), .C(rst_bF_buf39), .Y(_6746__10_) );
	OAI21X1 OAI21X1_3312 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf2), .B(_7320__bF_buf0), .C(csr_gpr_iu_csr_sscratch_11_), .Y(_7359_) );
	NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_7304__bF_buf6_bF_buf2), .Y(_7360_) );
	NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf0), .B(_7360_), .Y(_7361_) );
	AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_7359_), .B(_7361_), .C(rst_bF_buf38), .Y(_6746__11_) );
	OAI21X1 OAI21X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_12_), .Y(_7362_) );
	NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_7304__bF_buf4), .Y(_7363_) );
	NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf3), .B(_7363_), .Y(_7364_) );
	AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_7362_), .B(_7364_), .C(rst_bF_buf37), .Y(_6746__12_) );
	INVX1 INVX1_1225 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_13_), .Y(_7365_) );
	NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13_bF_buf3), .B(_7319__bF_buf3), .Y(_7366_) );
	OAI21X1 OAI21X1_3314 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_7366__bF_buf3), .C(_6879__bF_buf30), .Y(_7367_) );
	AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_7365_), .B(_7366__bF_buf2), .C(_7367_), .Y(_6746__13_) );
	OAI21X1 OAI21X1_3315 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_14_), .Y(_7368_) );
	INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .Y(_7369_) );
	NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7304__bF_buf2), .Y(_7370_) );
	NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf2), .B(_7370_), .Y(_7371_) );
	AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_7368_), .B(_7371_), .C(rst_bF_buf36), .Y(_6746__14_) );
	INVX1 INVX1_1226 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_15_), .Y(_7372_) );
	OAI21X1 OAI21X1_3316 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf0), .B(_7366__bF_buf1), .C(_6879__bF_buf29), .Y(_7373_) );
	AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_7372_), .B(_7366__bF_buf0), .C(_7373_), .Y(_6746__15_) );
	OAI21X1 OAI21X1_3317 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_7320__bF_buf1), .C(csr_gpr_iu_csr_sscratch_16_), .Y(_7374_) );
	INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .Y(_7375_) );
	NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_7304__bF_buf0), .Y(_7376_) );
	NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf1), .B(_7376_), .Y(_7377_) );
	AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_7374_), .B(_7377_), .C(rst_bF_buf35), .Y(_6746__16_) );
	INVX1 INVX1_1227 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_17_), .Y(_7378_) );
	OAI21X1 OAI21X1_3318 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf0), .B(_7366__bF_buf3), .C(_6879__bF_buf28), .Y(_7379_) );
	AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_7378_), .B(_7366__bF_buf2), .C(_7379_), .Y(_6746__17_) );
	OAI21X1 OAI21X1_3319 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf1), .B(_7320__bF_buf0), .C(csr_gpr_iu_csr_sscratch_18_), .Y(_7380_) );
	INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .Y(_7381_) );
	NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_7304__bF_buf13_bF_buf1), .Y(_7382_) );
	NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf0), .B(_7382_), .Y(_7383_) );
	AOI21X1 AOI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_7380_), .B(_7383_), .C(rst_bF_buf34), .Y(_6746__18_) );
	INVX1 INVX1_1228 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_19_), .Y(_7384_) );
	OAI21X1 OAI21X1_3320 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_7366__bF_buf1), .C(_6879__bF_buf27), .Y(_7385_) );
	AOI21X1 AOI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_7384_), .B(_7366__bF_buf0), .C(_7385_), .Y(_6746__19_) );
	OAI21X1 OAI21X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf1), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_20_), .Y(_7386_) );
	INVX1 INVX1_1229 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .Y(_7387_) );
	NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_7304__bF_buf11_bF_buf1), .Y(_7388_) );
	NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .B(_7388_), .Y(_7389_) );
	AOI21X1 AOI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_7386_), .B(_7389_), .C(rst_bF_buf33), .Y(_6746__20_) );
	INVX1 INVX1_1230 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_21_), .Y(_7390_) );
	OAI21X1 OAI21X1_3322 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_7366__bF_buf3), .C(_6879__bF_buf26), .Y(_7391_) );
	AOI21X1 AOI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_7390_), .B(_7366__bF_buf2), .C(_7391_), .Y(_6746__21_) );
	OAI21X1 OAI21X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf1), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_22_), .Y(_7392_) );
	INVX1 INVX1_1231 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .Y(_7393_) );
	NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7304__bF_buf9_bF_buf1), .Y(_7394_) );
	NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf3), .B(_7394_), .Y(_7395_) );
	AOI21X1 AOI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_7392_), .B(_7395_), .C(rst_bF_buf32), .Y(_6746__22_) );
	INVX1 INVX1_1232 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_23_), .Y(_7396_) );
	OAI21X1 OAI21X1_3324 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf3), .B(_7366__bF_buf1), .C(_6879__bF_buf25), .Y(_7397_) );
	AOI21X1 AOI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_7396_), .B(_7366__bF_buf0), .C(_7397_), .Y(_6746__23_) );
	OAI21X1 OAI21X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf1), .B(_7320__bF_buf1), .C(csr_gpr_iu_csr_sscratch_24_), .Y(_7398_) );
	INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .Y(_7399_) );
	NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_7399_), .B(_7304__bF_buf7_bF_buf1), .Y(_7400_) );
	NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf2), .B(_7400_), .Y(_7401_) );
	AOI21X1 AOI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_7398_), .B(_7401_), .C(rst_bF_buf31), .Y(_6746__24_) );
	INVX1 INVX1_1233 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_25_), .Y(_7402_) );
	OAI21X1 OAI21X1_3326 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_7366__bF_buf3), .C(_6879__bF_buf24), .Y(_7403_) );
	AOI21X1 AOI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_7402_), .B(_7366__bF_buf2), .C(_7403_), .Y(_6746__25_) );
	OAI21X1 OAI21X1_3327 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf1), .B(_7320__bF_buf0), .C(csr_gpr_iu_csr_sscratch_26_), .Y(_7404_) );
	INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .Y(_7405_) );
	NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7304__bF_buf5), .Y(_7406_) );
	NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf1), .B(_7406_), .Y(_7407_) );
	AOI21X1 AOI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_7404_), .B(_7407_), .C(rst_bF_buf30), .Y(_6746__26_) );
	INVX1 INVX1_1234 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_27_), .Y(_7408_) );
	OAI21X1 OAI21X1_3328 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_7366__bF_buf1), .C(_6879__bF_buf23), .Y(_7409_) );
	AOI21X1 AOI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_7408_), .B(_7366__bF_buf0), .C(_7409_), .Y(_6746__27_) );
	OAI21X1 OAI21X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_7320__bF_buf3), .C(csr_gpr_iu_csr_sscratch_28_), .Y(_7410_) );
	INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .Y(_7411_) );
	NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_7304__bF_buf3), .Y(_7412_) );
	NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf0), .B(_7412_), .Y(_7413_) );
	AOI21X1 AOI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_7410_), .B(_7413_), .C(rst_bF_buf29), .Y(_6746__28_) );
	INVX1 INVX1_1235 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_29_), .Y(_7414_) );
	OAI21X1 OAI21X1_3330 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_7366__bF_buf3), .C(_6879__bF_buf22), .Y(_7415_) );
	AOI21X1 AOI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_7414_), .B(_7366__bF_buf2), .C(_7415_), .Y(_6746__29_) );
	OAI21X1 OAI21X1_3331 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_7320__bF_buf2), .C(csr_gpr_iu_csr_sscratch_30_), .Y(_7416_) );
	NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_7304__bF_buf1), .Y(_7417_) );
	NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .B(_7417_), .Y(_7418_) );
	AOI21X1 AOI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_7416_), .B(_7418_), .C(rst_bF_buf28), .Y(_6746__30_) );
	INVX1 INVX1_1236 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_31_), .Y(_7419_) );
	OAI21X1 OAI21X1_3332 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf3), .B(_7366__bF_buf1), .C(_6879__bF_buf21), .Y(_7420_) );
	AOI21X1 AOI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_7419_), .B(_7366__bF_buf0), .C(_7420_), .Y(_6746__31_) );
	INVX1 INVX1_1237 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_0_), .Y(_7421_) );
	NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_2_), .Y(_7422_) );
	NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_7422_), .Y(_7423_) );
	INVX8 INVX8_62 ( .gnd(gnd), .vdd(vdd), .A(_7423_), .Y(_7424_) );
	INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .Y(_7425_) );
	NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf3), .B(_7425_), .Y(_7426_) );
	INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(_7426_), .Y(_7427_) );
	NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_7427_), .B(_7424__bF_buf3), .Y(_7428_) );
	INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_0_), .Y(_7429_) );
	NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_7303__bF_buf12_bF_buf3), .Y(_7430_) );
	NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf1), .B(_7310_), .Y(_7431_) );
	OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .B(biu_ins_20_bF_buf2), .Y(_7432_) );
	INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(_7432_), .Y(_7433_) );
	NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7433_), .Y(_7434_) );
	NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_7309__bF_buf2), .B(_7434__bF_buf4), .Y(_7435_) );
	AOI22X1 AOI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_7430_), .C(_7435__bF_buf6), .D(_7325_), .Y(_7436_) );
	INVX4 INVX4_17 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf5), .Y(_7437_) );
	OAI21X1 OAI21X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_7303__bF_buf11_bF_buf3), .C(_6879__bF_buf20), .Y(_7438_) );
	AOI21X1 AOI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_7437_), .B(_7303__bF_buf10_bF_buf3), .C(_7438_), .Y(_7439_) );
	OAI22X1 OAI22X1_647 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf27), .B(_7436_), .C(_7421_), .D(_7439__bF_buf4), .Y(_6739__0_) );
	INVX1 INVX1_1238 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_1_), .Y(_7440_) );
	INVX1 INVX1_1239 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .Y(_7441_) );
	NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_7441_), .B(_7303__bF_buf9_bF_buf3), .Y(_7442_) );
	AOI22X1 AOI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7442_), .C(_7435__bF_buf4), .D(_7329_), .Y(_7443_) );
	OAI22X1 OAI22X1_648 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf26), .B(_7443_), .C(_7440_), .D(_7439__bF_buf3), .Y(_6739__1_) );
	INVX1 INVX1_1240 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_2_), .Y(_7444_) );
	INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .Y(_7445_) );
	NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_7303__bF_buf8_bF_buf3), .Y(_7446_) );
	AOI22X1 AOI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7446_), .C(_7435__bF_buf3), .D(_7333_), .Y(_7447_) );
	OAI22X1 OAI22X1_649 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf25), .B(_7447_), .C(_7444_), .D(_7439__bF_buf2), .Y(_6739__2_) );
	INVX1 INVX1_1241 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_3_), .Y(_7448_) );
	INVX1 INVX1_1242 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_3_), .Y(_7449_) );
	NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_7303__bF_buf7_bF_buf3), .Y(_7450_) );
	AOI22X1 AOI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7450_), .C(_7435__bF_buf2), .D(_7336_), .Y(_7451_) );
	OAI22X1 OAI22X1_650 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf24), .B(_7451_), .C(_7448_), .D(_7439__bF_buf1), .Y(_6739__3_) );
	INVX1 INVX1_1243 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_4_), .Y(_7452_) );
	INVX1 INVX1_1244 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .Y(_7453_) );
	NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_7303__bF_buf6_bF_buf3), .Y(_7454_) );
	AOI22X1 AOI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_7454_), .C(_7435__bF_buf1), .D(_7339_), .Y(_7455_) );
	OAI22X1 OAI22X1_651 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf23), .B(_7455_), .C(_7452_), .D(_7439__bF_buf0), .Y(_6739__4_) );
	INVX1 INVX1_1245 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_5_), .Y(_7456_) );
	INVX1 INVX1_1246 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .Y(_7457_) );
	NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .B(_7303__bF_buf5_bF_buf3), .Y(_7458_) );
	AOI22X1 AOI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_7458_), .C(_7435__bF_buf0), .D(_7342_), .Y(_7459_) );
	OAI22X1 OAI22X1_652 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf22), .B(_7459_), .C(_7456_), .D(_7439__bF_buf4), .Y(_6739__5_) );
	INVX1 INVX1_1247 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_6_), .Y(_7460_) );
	INVX1 INVX1_1248 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .Y(_7461_) );
	NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_7303__bF_buf4_bF_buf3), .Y(_7462_) );
	AOI22X1 AOI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_7462_), .C(_7435__bF_buf6), .D(_7345_), .Y(_7463_) );
	OAI22X1 OAI22X1_653 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf21), .B(_7463_), .C(_7460_), .D(_7439__bF_buf3), .Y(_6739__6_) );
	INVX1 INVX1_1249 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_7_), .Y(_7464_) );
	INVX1 INVX1_1250 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .Y(_7465_) );
	NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .B(_7303__bF_buf3_bF_buf3), .Y(_7466_) );
	AOI22X1 AOI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_7466_), .C(_7435__bF_buf5), .D(_7348_), .Y(_7467_) );
	OAI22X1 OAI22X1_654 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf20), .B(_7467_), .C(_7464_), .D(_7439__bF_buf2), .Y(_6739__7_) );
	INVX1 INVX1_1251 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_8_), .Y(_7468_) );
	INVX1 INVX1_1252 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .Y(_7469_) );
	NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_7469_), .B(_7303__bF_buf2), .Y(_7470_) );
	AOI22X1 AOI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_7470_), .C(_7435__bF_buf4), .D(_7351_), .Y(_7471_) );
	OAI22X1 OAI22X1_655 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf19), .B(_7471_), .C(_7468_), .D(_7439__bF_buf1), .Y(_6739__8_) );
	INVX1 INVX1_1253 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_9_), .Y(_7472_) );
	INVX1 INVX1_1254 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .Y(_7473_) );
	NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7303__bF_buf1), .Y(_7474_) );
	AOI22X1 AOI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_7474_), .C(_7435__bF_buf3), .D(_7354_), .Y(_7475_) );
	OAI22X1 OAI22X1_656 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf18), .B(_7475_), .C(_7472_), .D(_7439__bF_buf0), .Y(_6739__9_) );
	INVX1 INVX1_1255 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_10_), .Y(_7476_) );
	INVX1 INVX1_1256 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .Y(_7477_) );
	NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_7477_), .B(_7303__bF_buf0), .Y(_7478_) );
	AOI22X1 AOI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7478_), .C(_7435__bF_buf2), .D(_7357_), .Y(_7479_) );
	OAI22X1 OAI22X1_657 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf17), .B(_7479_), .C(_7476_), .D(_7439__bF_buf4), .Y(_6739__10_) );
	INVX1 INVX1_1257 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_11_), .Y(_7480_) );
	INVX1 INVX1_1258 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .Y(_7481_) );
	NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .B(_7303__bF_buf14_bF_buf2), .Y(_7482_) );
	AOI22X1 AOI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7482_), .C(_7435__bF_buf1), .D(_7360_), .Y(_7483_) );
	OAI22X1 OAI22X1_658 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf16), .B(_7483_), .C(_7480_), .D(_7439__bF_buf3), .Y(_6739__11_) );
	INVX1 INVX1_1259 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_12_), .Y(_7484_) );
	INVX1 INVX1_1260 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .Y(_7485_) );
	NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_7303__bF_buf13_bF_buf2), .Y(_7486_) );
	AOI22X1 AOI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7486_), .C(_7435__bF_buf0), .D(_7363_), .Y(_7487_) );
	OAI22X1 OAI22X1_659 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf15), .B(_7487_), .C(_7484_), .D(_7439__bF_buf2), .Y(_6739__12_) );
	INVX1 INVX1_1261 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_13_), .Y(_7488_) );
	INVX1 INVX1_1262 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .Y(_7489_) );
	NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_7303__bF_buf12_bF_buf2), .Y(_7490_) );
	INVX1 INVX1_1263 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf2), .Y(_7491_) );
	NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_7491_), .B(_7304__bF_buf0), .Y(_7492_) );
	AOI22X1 AOI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_7490_), .B(_7428__bF_buf3), .C(_7435__bF_buf6), .D(_7492_), .Y(_7493_) );
	OAI22X1 OAI22X1_660 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf14), .B(_7493_), .C(_7488_), .D(_7439__bF_buf1), .Y(_6739__13_) );
	INVX1 INVX1_1264 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_14_), .Y(_7494_) );
	INVX1 INVX1_1265 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .Y(_7495_) );
	NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_7495_), .B(_7303__bF_buf11_bF_buf2), .Y(_7496_) );
	AOI22X1 AOI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_7496_), .C(_7435__bF_buf5), .D(_7370_), .Y(_7497_) );
	OAI22X1 OAI22X1_661 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf13), .B(_7497_), .C(_7494_), .D(_7439__bF_buf0), .Y(_6739__14_) );
	INVX1 INVX1_1266 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_15_), .Y(_7498_) );
	INVX1 INVX1_1267 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .Y(_7499_) );
	NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_7303__bF_buf10_bF_buf2), .Y(_7500_) );
	NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_6978_), .B(_7304__bF_buf14_bF_buf0), .Y(_7501_) );
	AOI22X1 AOI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_7500_), .B(_7428__bF_buf1), .C(_7435__bF_buf4), .D(_7501_), .Y(_7502_) );
	OAI22X1 OAI22X1_662 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf12), .B(_7502_), .C(_7498_), .D(_7439__bF_buf4), .Y(_6739__15_) );
	INVX1 INVX1_1268 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_16_), .Y(_7503_) );
	INVX1 INVX1_1269 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .Y(_7504_) );
	NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .B(_7303__bF_buf9_bF_buf2), .Y(_7505_) );
	AOI22X1 AOI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_7505_), .C(_7435__bF_buf3), .D(_7376_), .Y(_7506_) );
	OAI22X1 OAI22X1_663 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf11), .B(_7506_), .C(_7503_), .D(_7439__bF_buf3), .Y(_6739__16_) );
	INVX1 INVX1_1270 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_17_), .Y(_7507_) );
	INVX1 INVX1_1271 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .Y(_7508_) );
	NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7303__bF_buf8_bF_buf2), .Y(_7509_) );
	NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_7304__bF_buf13_bF_buf0), .Y(_7510_) );
	AOI22X1 AOI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(_7509_), .B(_7428__bF_buf8), .C(_7435__bF_buf2), .D(_7510_), .Y(_7511_) );
	OAI22X1 OAI22X1_664 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf10), .B(_7511_), .C(_7507_), .D(_7439__bF_buf2), .Y(_6739__17_) );
	INVX1 INVX1_1272 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_18_), .Y(_7512_) );
	INVX1 INVX1_1273 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .Y(_7513_) );
	NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_7513_), .B(_7303__bF_buf7_bF_buf2), .Y(_7514_) );
	AOI22X1 AOI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_7514_), .C(_7435__bF_buf1), .D(_7382_), .Y(_7515_) );
	OAI22X1 OAI22X1_665 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf9), .B(_7515_), .C(_7512_), .D(_7439__bF_buf1), .Y(_6739__18_) );
	INVX1 INVX1_1274 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_19_), .Y(_7516_) );
	INVX1 INVX1_1275 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .Y(_7517_) );
	NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_7517_), .B(_7303__bF_buf6_bF_buf2), .Y(_7518_) );
	AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5_bF_buf2), .B(addr_csr_19_bF_buf2), .Y(_7519_) );
	AOI22X1 AOI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7518_), .C(_7519_), .D(_7435__bF_buf0), .Y(_7520_) );
	OAI22X1 OAI22X1_666 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf8), .B(_7520_), .C(_7516_), .D(_7439__bF_buf0), .Y(_6739__19_) );
	INVX1 INVX1_1276 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_20_), .Y(_7521_) );
	INVX1 INVX1_1277 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .Y(_7522_) );
	NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_7522_), .B(_7303__bF_buf4_bF_buf2), .Y(_7523_) );
	AOI22X1 AOI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7523_), .C(_7435__bF_buf6), .D(_7388_), .Y(_7524_) );
	OAI22X1 OAI22X1_667 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf7), .B(_7524_), .C(_7521_), .D(_7439__bF_buf4), .Y(_6739__20_) );
	INVX1 INVX1_1278 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_21_), .Y(_7525_) );
	INVX1 INVX1_1279 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .Y(_7526_) );
	NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_7526_), .B(_7303__bF_buf3_bF_buf2), .Y(_7527_) );
	AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf2), .B(addr_csr_21_bF_buf2), .Y(_7528_) );
	AOI22X1 AOI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7527_), .C(_7528_), .D(_7435__bF_buf5), .Y(_7529_) );
	OAI22X1 OAI22X1_668 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf6), .B(_7529_), .C(_7525_), .D(_7439__bF_buf3), .Y(_6739__21_) );
	INVX1 INVX1_1280 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_22_), .Y(_7530_) );
	INVX1 INVX1_1281 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .Y(_7531_) );
	NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_7531_), .B(_7303__bF_buf1), .Y(_7532_) );
	AOI22X1 AOI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_7532_), .C(_7435__bF_buf4), .D(_7394_), .Y(_7533_) );
	OAI22X1 OAI22X1_669 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .B(_7533_), .C(_7530_), .D(_7439__bF_buf2), .Y(_6739__22_) );
	INVX1 INVX1_1282 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_23_), .Y(_7534_) );
	INVX1 INVX1_1283 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .Y(_7535_) );
	NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_7535_), .B(_7303__bF_buf0), .Y(_7536_) );
	NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_7304__bF_buf12_bF_buf0), .Y(_7537_) );
	AOI22X1 AOI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(_7536_), .B(_7428__bF_buf2), .C(_7435__bF_buf3), .D(_7537_), .Y(_7538_) );
	OAI22X1 OAI22X1_670 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_7538_), .C(_7534_), .D(_7439__bF_buf1), .Y(_6739__23_) );
	INVX1 INVX1_1284 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_24_), .Y(_7539_) );
	INVX1 INVX1_1285 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .Y(_7540_) );
	NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .B(_7303__bF_buf14_bF_buf1), .Y(_7541_) );
	AOI22X1 AOI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_7541_), .C(_7435__bF_buf2), .D(_7400_), .Y(_7542_) );
	OAI22X1 OAI22X1_671 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_7542_), .C(_7539_), .D(_7439__bF_buf0), .Y(_6739__24_) );
	INVX1 INVX1_1286 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_25_), .Y(_7543_) );
	INVX1 INVX1_1287 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .Y(_7544_) );
	NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_7544_), .B(_7303__bF_buf13_bF_buf1), .Y(_7545_) );
	AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12_bF_buf1), .B(addr_csr_25_bF_buf2), .Y(_7546_) );
	AOI22X1 AOI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_7545_), .C(_7546_), .D(_7435__bF_buf1), .Y(_7547_) );
	OAI22X1 OAI22X1_672 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_7547_), .C(_7543_), .D(_7439__bF_buf4), .Y(_6739__25_) );
	INVX1 INVX1_1288 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_26_), .Y(_7548_) );
	INVX1 INVX1_1289 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .Y(_7549_) );
	NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_7549_), .B(_7303__bF_buf11_bF_buf1), .Y(_7550_) );
	AOI22X1 AOI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_7550_), .C(_7435__bF_buf0), .D(_7406_), .Y(_7551_) );
	OAI22X1 OAI22X1_673 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_7551_), .C(_7548_), .D(_7439__bF_buf3), .Y(_6739__26_) );
	INVX1 INVX1_1290 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_27_), .Y(_7552_) );
	INVX1 INVX1_1291 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_27_), .Y(_7553_) );
	NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_7553_), .B(_7303__bF_buf10_bF_buf1), .Y(_7554_) );
	INVX1 INVX1_1292 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf2), .Y(_7555_) );
	NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_7555_), .B(_7304__bF_buf11_bF_buf0), .Y(_7556_) );
	AOI22X1 AOI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(_7554_), .B(_7428__bF_buf7), .C(_7435__bF_buf6), .D(_7556_), .Y(_7557_) );
	OAI22X1 OAI22X1_674 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_7557_), .C(_7552_), .D(_7439__bF_buf2), .Y(_6739__27_) );
	INVX1 INVX1_1293 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_28_), .Y(_7558_) );
	INVX1 INVX1_1294 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .Y(_7559_) );
	NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_7559_), .B(_7303__bF_buf9_bF_buf1), .Y(_7560_) );
	AOI22X1 AOI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7560_), .C(_7435__bF_buf5), .D(_7412_), .Y(_7561_) );
	OAI22X1 OAI22X1_675 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf70), .B(_7561_), .C(_7558_), .D(_7439__bF_buf1), .Y(_6739__28_) );
	INVX1 INVX1_1295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_29_), .Y(_7562_) );
	INVX1 INVX1_1296 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .Y(_7563_) );
	NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .B(_7303__bF_buf8_bF_buf1), .Y(_7564_) );
	AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7_bF_buf1), .B(addr_csr_29_bF_buf2), .Y(_7565_) );
	AOI22X1 AOI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7564_), .C(_7565_), .D(_7435__bF_buf4), .Y(_7566_) );
	OAI22X1 OAI22X1_676 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf69), .B(_7566_), .C(_7562_), .D(_7439__bF_buf0), .Y(_6739__29_) );
	INVX1 INVX1_1297 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_30_), .Y(_7567_) );
	INVX1 INVX1_1298 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .Y(_7568_) );
	NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_7568_), .B(_7303__bF_buf6_bF_buf1), .Y(_7569_) );
	AOI22X1 AOI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7569_), .C(_7435__bF_buf3), .D(_7417_), .Y(_7570_) );
	OAI22X1 OAI22X1_677 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_7570_), .C(_7567_), .D(_7439__bF_buf4), .Y(_6739__30_) );
	INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf3), .Y(_7571_) );
	INVX1 INVX1_1299 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .Y(_7572_) );
	NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_7572_), .B(_7303__bF_buf5_bF_buf1), .Y(_7573_) );
	NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_7278_), .B(_7304__bF_buf10_bF_buf0), .Y(_7574_) );
	AOI22X1 AOI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(_7573_), .B(_7428__bF_buf3), .C(_7435__bF_buf2), .D(_7574_), .Y(_7575_) );
	OAI22X1 OAI22X1_678 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf67), .B(_7575_), .C(_7571_), .D(_7439__bF_buf3), .Y(_6739__31_) );
	INVX1 INVX1_1300 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_0_), .Y(_7576_) );
	INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .Y(_7577_) );
	NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7303__bF_buf4_bF_buf1), .Y(_7578_) );
	INVX1 INVX1_1301 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf1), .Y(_7579_) );
	NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf0), .B(_7579_), .Y(_7580_) );
	NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_7310_), .B(_7580_), .Y(_7581_) );
	INVX1 INVX1_1302 ( .gnd(gnd), .vdd(vdd), .A(_7581_), .Y(_7582_) );
	NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7582_), .Y(_7583_) );
	NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf3), .B(_7309__bF_buf1), .Y(_7584_) );
	AOI22X1 AOI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_7578_), .C(_7584__bF_buf5), .D(_7325_), .Y(_7585_) );
	INVX8 INVX8_63 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf4), .Y(_7586_) );
	AOI21X1 AOI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_7586__bF_buf5), .B(_7303__bF_buf3_bF_buf1), .C(_7438_), .Y(_7587_) );
	OAI22X1 OAI22X1_679 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf66), .B(_7585_), .C(_7576_), .D(_7587_), .Y(_6742__0_) );
	INVX1 INVX1_1303 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_1_), .Y(_7588_) );
	INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .Y(_7589_) );
	NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_7303__bF_buf2), .Y(_7590_) );
	AOI22X1 AOI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_7590_), .C(_7584__bF_buf3), .D(_7329_), .Y(_7591_) );
	OAI22X1 OAI22X1_680 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf65), .B(_7591_), .C(_7588_), .D(_7587_), .Y(_6742__1_) );
	OAI21X1 OAI21X1_3334 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf2), .B(_7309__bF_buf0), .C(csr_gpr_iu_csr_sepc_2_), .Y(_7592_) );
	OAI21X1 OAI21X1_3335 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7586__bF_buf4), .C(_7592_), .Y(_7593_) );
	INVX8 INVX8_64 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .Y(_7594_) );
	INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .Y(_7595_) );
	OAI21X1 OAI21X1_3336 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .B(csr_gpr_iu_cause_3_), .C(_7445_), .Y(_7596_) );
	OAI21X1 OAI21X1_3337 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_0_), .B(_7441_), .C(_7453_), .Y(_7597_) );
	NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_7596_), .B(_7597_), .Y(_7598_) );
	NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .B(csr_gpr_iu_cause_31_bF_buf6), .Y(_7599_) );
	NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7522_), .C(_7599_), .Y(_7600_) );
	NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .B(csr_gpr_iu_cause_31_bF_buf4), .Y(_7601_) );
	NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_7504_), .C(_7601_), .Y(_7602_) );
	NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_7600_), .B(_7602_), .Y(_7603_) );
	NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_7603_), .Y(_7604_) );
	NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .B(csr_gpr_iu_cause_27_), .Y(_7605_) );
	NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .B(csr_gpr_iu_cause_31_bF_buf1), .Y(_7606_) );
	NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .B(csr_gpr_iu_cause_31_bF_buf6), .Y(_7607_) );
	NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_7605_), .B(_7606_), .C(_7607_), .Y(_7608_) );
	NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .B(csr_gpr_iu_cause_31_bF_buf4), .Y(_7609_) );
	NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .B(csr_gpr_iu_cause_31_bF_buf2), .Y(_7610_) );
	NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_7568_), .B(_7609_), .C(_7610_), .Y(_7611_) );
	NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_7611_), .B(_7608_), .Y(_7612_) );
	NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .B(csr_gpr_iu_cause_31_bF_buf0), .Y(_7613_) );
	NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7485_), .C(_7613_), .Y(_7614_) );
	NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .B(csr_gpr_iu_cause_31_bF_buf5), .Y(_7615_) );
	NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .B(_7615_), .Y(_7616_) );
	NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_7616_), .B(_7614_), .Y(_7617_) );
	AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .B(_7469_), .Y(_7618_) );
	NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_7618_), .Y(_7619_) );
	NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_7619_), .Y(_7620_) );
	XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_7620_), .B(_7595_), .Y(_7621_) );
	INVX1 INVX1_1304 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .Y(_7622_) );
	AOI21X1 AOI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(csr_gpr_iu_csr_sepc_2_), .C(_7303__bF_buf1), .Y(_7623_) );
	OAI21X1 OAI21X1_3338 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7622_), .C(_7623_), .Y(_7624_) );
	OAI21X1 OAI21X1_3339 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf0), .B(_7593_), .C(_7624_), .Y(_7625_) );
	NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf64), .B(csr_gpr_iu_csr_sepc_2_), .Y(_7626_) );
	OAI21X1 OAI21X1_3340 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf63), .B(_7625_), .C(_7626_), .Y(_6742__2_) );
	OAI21X1 OAI21X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf1), .B(_7309__bF_buf3), .C(csr_gpr_iu_csr_sepc_3_), .Y(_7627_) );
	OAI21X1 OAI21X1_3342 ( .gnd(gnd), .vdd(vdd), .A(_6895_), .B(_7586__bF_buf3), .C(_7627_), .Y(_7628_) );
	INVX1 INVX1_1305 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .Y(_7629_) );
	INVX1 INVX1_1306 ( .gnd(gnd), .vdd(vdd), .A(_7620_), .Y(_7630_) );
	OAI21X1 OAI21X1_3343 ( .gnd(gnd), .vdd(vdd), .A(_7595_), .B(_7630_), .C(_7629_), .Y(_7631_) );
	INVX1 INVX1_1307 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .Y(_7632_) );
	NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_7603_), .C(_7618_), .Y(_7633_) );
	NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_7632_), .B(_7633_), .Y(_7634_) );
	NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(biu_pc_3_), .C(_7634_), .Y(_7635_) );
	NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_7635_), .B(_7631_), .Y(_7636_) );
	INVX1 INVX1_1308 ( .gnd(gnd), .vdd(vdd), .A(_7636_), .Y(_7637_) );
	NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7637_), .Y(_7638_) );
	NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_3_), .B(_7428__bF_buf8), .Y(_7639_) );
	OAI21X1 OAI21X1_3344 ( .gnd(gnd), .vdd(vdd), .A(_7639_), .B(_7638_), .C(_7304__bF_buf8_bF_buf0), .Y(_7640_) );
	OAI21X1 OAI21X1_3345 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf0), .B(_7628_), .C(_7640_), .Y(_7641_) );
	NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf62), .B(csr_gpr_iu_csr_sepc_3_), .Y(_7642_) );
	OAI21X1 OAI21X1_3346 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf61), .B(_7641_), .C(_7642_), .Y(_6742__3_) );
	OAI21X1 OAI21X1_3347 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf0), .B(_7309__bF_buf2), .C(csr_gpr_iu_csr_sepc_4_), .Y(_7643_) );
	OAI21X1 OAI21X1_3348 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_7586__bF_buf2), .C(_7643_), .Y(_7644_) );
	INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .Y(_7645_) );
	XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_7635_), .B(_7645_), .Y(_7646_) );
	INVX1 INVX1_1309 ( .gnd(gnd), .vdd(vdd), .A(_7646_), .Y(_7647_) );
	NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7647_), .Y(_7648_) );
	NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_4_), .B(_7428__bF_buf7), .Y(_7649_) );
	OAI21X1 OAI21X1_3349 ( .gnd(gnd), .vdd(vdd), .A(_7649_), .B(_7648_), .C(_7304__bF_buf6_bF_buf0), .Y(_7650_) );
	OAI21X1 OAI21X1_3350 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_7644_), .C(_7650_), .Y(_7651_) );
	NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf60), .B(csr_gpr_iu_csr_sepc_4_), .Y(_7652_) );
	OAI21X1 OAI21X1_3351 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf59), .B(_7651_), .C(_7652_), .Y(_6742__4_) );
	INVX1 INVX1_1310 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_5_), .Y(_7653_) );
	NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_7645_), .B(_7635_), .Y(_7654_) );
	NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .B(_7654_), .Y(_7655_) );
	INVX1 INVX1_1311 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .Y(_7656_) );
	OAI21X1 OAI21X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_7645_), .B(_7635_), .C(_7656_), .Y(_7657_) );
	AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .B(_7657_), .Y(_7658_) );
	AOI21X1 AOI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7653_), .C(_7303__bF_buf0), .Y(_7659_) );
	OAI21X1 OAI21X1_3353 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7658_), .C(_7659_), .Y(_7660_) );
	OAI21X1 OAI21X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf3), .B(_7309__bF_buf1), .C(csr_gpr_iu_csr_sepc_5_), .Y(_7661_) );
	OAI21X1 OAI21X1_3355 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_7586__bF_buf1), .C(_7661_), .Y(_7662_) );
	AOI21X1 AOI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(_7303__bF_buf14_bF_buf0), .C(rst_bF_buf58), .Y(_7663_) );
	AOI22X1 AOI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf57), .B(_7653_), .C(_7663_), .D(_7660_), .Y(_6742__5_) );
	OAI21X1 OAI21X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf2), .B(_7309__bF_buf0), .C(csr_gpr_iu_csr_sepc_6_), .Y(_7664_) );
	OAI21X1 OAI21X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_7586__bF_buf0), .C(_7664_), .Y(_7665_) );
	INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .Y(_7666_) );
	XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .B(_7666_), .Y(_7667_) );
	AOI21X1 AOI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(csr_gpr_iu_csr_sepc_6_), .C(_7303__bF_buf13_bF_buf0), .Y(_7668_) );
	OAI21X1 OAI21X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7667_), .C(_7668_), .Y(_7669_) );
	OAI21X1 OAI21X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_7665_), .C(_7669_), .Y(_7670_) );
	NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf56), .B(csr_gpr_iu_csr_sepc_6_), .Y(_7671_) );
	OAI21X1 OAI21X1_3360 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf55), .B(_7670_), .C(_7671_), .Y(_6742__6_) );
	INVX1 INVX1_1312 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_7_), .Y(_7672_) );
	INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .Y(_7673_) );
	OAI21X1 OAI21X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_7666_), .B(_7655_), .C(_7673_), .Y(_7674_) );
	NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_7666_), .B(_7655_), .Y(_7675_) );
	NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .B(_7675_), .Y(_7676_) );
	AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_7676_), .B(_7674_), .Y(_7677_) );
	AOI21X1 AOI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7672_), .C(_7303__bF_buf12_bF_buf0), .Y(_7678_) );
	OAI21X1 OAI21X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7677_), .C(_7678_), .Y(_7679_) );
	OAI21X1 OAI21X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf1), .B(_7309__bF_buf3), .C(csr_gpr_iu_csr_sepc_7_), .Y(_7680_) );
	OAI21X1 OAI21X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_7586__bF_buf5), .C(_7680_), .Y(_7681_) );
	AOI21X1 AOI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_7681_), .B(_7303__bF_buf11_bF_buf0), .C(rst_bF_buf54), .Y(_7682_) );
	AOI22X1 AOI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf53), .B(_7672_), .C(_7682_), .D(_7679_), .Y(_6742__7_) );
	INVX1 INVX1_1313 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_8_), .Y(_7683_) );
	NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(biu_pc_3_), .Y(_7684_) );
	NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .B(biu_pc_5_), .Y(_7685_) );
	NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_7684_), .B(_7685_), .Y(_7686_) );
	NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .B(_7686_), .Y(_7687_) );
	NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(_7687_), .Y(_7688_) );
	NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_7688_), .B(_7620_), .Y(_7689_) );
	XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_7689_), .B(biu_pc_8_), .Y(_7690_) );
	AOI21X1 AOI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7683_), .C(_7303__bF_buf10_bF_buf0), .Y(_7691_) );
	OAI21X1 OAI21X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7690_), .C(_7691_), .Y(_7692_) );
	NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_7586__bF_buf4), .Y(_7693_) );
	OAI21X1 OAI21X1_3366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_8_), .B(_7584__bF_buf2), .C(_7303__bF_buf9_bF_buf0), .Y(_7694_) );
	OAI21X1 OAI21X1_3367 ( .gnd(gnd), .vdd(vdd), .A(_7693_), .B(_7694_), .C(_7692_), .Y(_7695_) );
	NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf19), .B(_7695_), .Y(_7696_) );
	OAI21X1 OAI21X1_3368 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf18), .B(_7683_), .C(_7696_), .Y(_6742__8_) );
	INVX1 INVX1_1314 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_9_), .Y(_7697_) );
	INVX1 INVX1_1315 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .Y(_7698_) );
	INVX1 INVX1_1316 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .Y(_7699_) );
	NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_7699_), .B(_7689_), .Y(_7700_) );
	XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_7700_), .B(_7698_), .Y(_7701_) );
	AOI21X1 AOI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7697_), .C(_7303__bF_buf8_bF_buf0), .Y(_7702_) );
	OAI21X1 OAI21X1_3369 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(_7701_), .C(_7702_), .Y(_7703_) );
	NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_7586__bF_buf3), .Y(_7704_) );
	OAI21X1 OAI21X1_3370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_9_), .B(_7584__bF_buf1), .C(_7303__bF_buf7_bF_buf0), .Y(_7705_) );
	OAI21X1 OAI21X1_3371 ( .gnd(gnd), .vdd(vdd), .A(_7704_), .B(_7705_), .C(_7703_), .Y(_7706_) );
	NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf17), .B(_7706_), .Y(_7707_) );
	OAI21X1 OAI21X1_3372 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf16), .B(_7697_), .C(_7707_), .Y(_6742__9_) );
	INVX1 INVX1_1317 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_10_), .Y(_7708_) );
	INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .Y(_7709_) );
	NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .B(biu_pc_9_), .Y(_7710_) );
	OAI21X1 OAI21X1_3373 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7676_), .C(_7709_), .Y(_7711_) );
	NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .B(biu_pc_9_), .C(_7688_), .Y(_7712_) );
	NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_7709_), .B(_7712_), .Y(_7713_) );
	NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .B(_7620_), .Y(_7714_) );
	AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_7711_), .B(_7714_), .Y(_7715_) );
	AOI21X1 AOI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7708_), .C(_7303__bF_buf6_bF_buf0), .Y(_7716_) );
	OAI21X1 OAI21X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7715_), .C(_7716_), .Y(_7717_) );
	OAI21X1 OAI21X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf0), .B(_7309__bF_buf2), .C(csr_gpr_iu_csr_sepc_10_), .Y(_7718_) );
	OAI21X1 OAI21X1_3376 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_7586__bF_buf2), .C(_7718_), .Y(_7719_) );
	AOI21X1 AOI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_7719_), .B(_7303__bF_buf5_bF_buf0), .C(rst_bF_buf52), .Y(_7720_) );
	AOI22X1 AOI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf51), .B(_7708_), .C(_7720_), .D(_7717_), .Y(_6742__10_) );
	OAI21X1 OAI21X1_3377 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf3), .B(_7309__bF_buf1), .C(csr_gpr_iu_csr_sepc_11_), .Y(_7721_) );
	OAI21X1 OAI21X1_3378 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_7586__bF_buf1), .C(_7721_), .Y(_7722_) );
	INVX1 INVX1_1318 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .Y(_7723_) );
	NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_7723_), .B(_7714_), .Y(_7724_) );
	INVX1 INVX1_1319 ( .gnd(gnd), .vdd(vdd), .A(_7714_), .Y(_7725_) );
	NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(_7725_), .Y(_7726_) );
	AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_7726_), .B(_7724_), .Y(_7727_) );
	INVX1 INVX1_1320 ( .gnd(gnd), .vdd(vdd), .A(_7727_), .Y(_7728_) );
	AOI21X1 AOI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(csr_gpr_iu_csr_sepc_11_), .C(_7303__bF_buf4_bF_buf0), .Y(_7729_) );
	OAI21X1 OAI21X1_3379 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7728_), .C(_7729_), .Y(_7730_) );
	OAI21X1 OAI21X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_7722_), .C(_7730_), .Y(_7731_) );
	NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf50), .B(csr_gpr_iu_csr_sepc_11_), .Y(_7732_) );
	OAI21X1 OAI21X1_3381 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf49), .B(_7731_), .C(_7732_), .Y(_6742__11_) );
	INVX1 INVX1_1321 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_12_), .Y(_7733_) );
	XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_7726_), .B(biu_pc_12_), .Y(_7734_) );
	AOI21X1 AOI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7733_), .C(_7303__bF_buf3_bF_buf0), .Y(_7735_) );
	OAI21X1 OAI21X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7734_), .C(_7735_), .Y(_7736_) );
	NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_7586__bF_buf0), .Y(_7737_) );
	OAI21X1 OAI21X1_3383 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_12_), .B(_7584__bF_buf0), .C(_7303__bF_buf2), .Y(_7738_) );
	OAI21X1 OAI21X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_7737_), .B(_7738_), .C(_7736_), .Y(_7739_) );
	NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf15), .B(_7739_), .Y(_7740_) );
	OAI21X1 OAI21X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf14), .B(_7733_), .C(_7740_), .Y(_6742__12_) );
	INVX1 INVX1_1322 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .Y(_7741_) );
	INVX1 INVX1_1323 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .Y(_7742_) );
	OAI21X1 OAI21X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(_7726_), .C(_7742_), .Y(_7743_) );
	INVX1 INVX1_1324 ( .gnd(gnd), .vdd(vdd), .A(_7743_), .Y(_7744_) );
	NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(biu_pc_12_), .C(biu_pc_13_), .Y(_7745_) );
	NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_7745_), .B(_7714_), .Y(_7746_) );
	OAI21X1 OAI21X1_3387 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_7744_), .C(_7428__bF_buf6), .Y(_7747_) );
	INVX1 INVX1_1325 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_13_), .Y(_7748_) );
	AOI21X1 AOI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(_7748_), .C(_7303__bF_buf1), .Y(_7749_) );
	OAI21X1 OAI21X1_3388 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf2), .B(_7309__bF_buf0), .C(csr_gpr_iu_csr_sepc_13_), .Y(_7750_) );
	OAI21X1 OAI21X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_7491_), .B(_7586__bF_buf5), .C(_7750_), .Y(_7751_) );
	AOI22X1 AOI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf0), .B(_7751_), .C(_7749_), .D(_7747_), .Y(_7752_) );
	NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf48), .B(csr_gpr_iu_csr_sepc_13_), .Y(_7753_) );
	OAI21X1 OAI21X1_3390 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf47), .B(_7752_), .C(_7753_), .Y(_6742__13_) );
	NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(_7746_), .Y(_7754_) );
	INVX1 INVX1_1326 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .Y(_7755_) );
	INVX1 INVX1_1327 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .Y(_7756_) );
	NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_7755_), .B(_7756_), .Y(_7757_) );
	OAI21X1 OAI21X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .B(_7757_), .C(_7428__bF_buf5), .Y(_7758_) );
	OAI21X1 OAI21X1_3392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_14_), .B(_7428__bF_buf4), .C(_7758_), .Y(_7759_) );
	OAI21X1 OAI21X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf4), .C(_7759_), .Y(_7760_) );
	AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_7586__bF_buf4), .B(csr_gpr_iu_csr_sepc_14_), .Y(_7761_) );
	OAI21X1 OAI21X1_3394 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7586__bF_buf3), .C(_7303__bF_buf14_bF_buf3), .Y(_7762_) );
	OAI21X1 OAI21X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_7761_), .B(_7762_), .C(_7760_), .Y(_7763_) );
	NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf46), .B(csr_gpr_iu_csr_sepc_14_), .Y(_7764_) );
	OAI21X1 OAI21X1_3396 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf45), .B(_7763_), .C(_7764_), .Y(_6742__14_) );
	INVX1 INVX1_1328 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_15_), .Y(_7765_) );
	INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .Y(_7766_) );
	XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_7757_), .B(_7766_), .Y(_7767_) );
	AOI21X1 AOI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7765_), .C(_7303__bF_buf13_bF_buf3), .Y(_7768_) );
	OAI21X1 OAI21X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7767_), .C(_7768_), .Y(_7769_) );
	NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf3), .B(_7586__bF_buf2), .Y(_7770_) );
	OAI21X1 OAI21X1_3398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_15_), .B(_7584__bF_buf5), .C(_7303__bF_buf12_bF_buf3), .Y(_7771_) );
	OAI21X1 OAI21X1_3399 ( .gnd(gnd), .vdd(vdd), .A(_7770_), .B(_7771_), .C(_7769_), .Y(_7772_) );
	NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf13), .B(_7772_), .Y(_7773_) );
	OAI21X1 OAI21X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf12), .B(_7765_), .C(_7773_), .Y(_6742__15_) );
	AOI21X1 AOI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_7757_), .B(biu_pc_15_), .C(biu_pc_16_), .Y(_7774_) );
	NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(biu_pc_15_), .Y(_7775_) );
	INVX1 INVX1_1329 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .Y(_7776_) );
	NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .B(_7776_), .Y(_7777_) );
	NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .B(_7756_), .Y(_7778_) );
	OAI21X1 OAI21X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_7778_), .B(_7774_), .C(_7428__bF_buf3), .Y(_7779_) );
	INVX1 INVX1_1330 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_16_), .Y(_7780_) );
	AOI21X1 AOI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7780_), .C(_7303__bF_buf11_bF_buf3), .Y(_7781_) );
	OAI21X1 OAI21X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf1), .B(_7309__bF_buf3), .C(csr_gpr_iu_csr_sepc_16_), .Y(_7782_) );
	OAI21X1 OAI21X1_3403 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_7586__bF_buf1), .C(_7782_), .Y(_7783_) );
	AOI22X1 AOI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf3), .B(_7783_), .C(_7781_), .D(_7779_), .Y(_7784_) );
	NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf44), .B(csr_gpr_iu_csr_sepc_16_), .Y(_7785_) );
	OAI21X1 OAI21X1_3404 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf43), .B(_7784_), .C(_7785_), .Y(_6742__16_) );
	NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(_7778_), .Y(_7786_) );
	INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .Y(_7787_) );
	NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .B(_7745_), .Y(_7788_) );
	AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_7788_), .B(biu_pc_16_), .Y(_7789_) );
	NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_7789_), .B(_7725_), .Y(_7790_) );
	NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .B(_7790_), .Y(_7791_) );
	OAI21X1 OAI21X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_7786_), .C(_7428__bF_buf2), .Y(_7792_) );
	INVX1 INVX1_1331 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_17_), .Y(_7793_) );
	AOI21X1 AOI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7793_), .C(_7303__bF_buf9_bF_buf3), .Y(_7794_) );
	OAI21X1 OAI21X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf0), .B(_7309__bF_buf2), .C(csr_gpr_iu_csr_sepc_17_), .Y(_7795_) );
	OAI21X1 OAI21X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_7586__bF_buf0), .C(_7795_), .Y(_7796_) );
	AOI22X1 AOI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8_bF_buf3), .B(_7796_), .C(_7794_), .D(_7792_), .Y(_7797_) );
	NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf42), .B(csr_gpr_iu_csr_sepc_17_), .Y(_7798_) );
	OAI21X1 OAI21X1_3408 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf41), .B(_7797_), .C(_7798_), .Y(_6742__17_) );
	INVX1 INVX1_1332 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_18_), .Y(_7799_) );
	INVX1 INVX1_1333 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .Y(_7800_) );
	XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_7800_), .Y(_7801_) );
	AOI21X1 AOI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7799_), .C(_7303__bF_buf7_bF_buf3), .Y(_7802_) );
	OAI21X1 OAI21X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7801_), .C(_7802_), .Y(_7803_) );
	NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_7586__bF_buf5), .Y(_7804_) );
	OAI21X1 OAI21X1_3410 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_18_), .B(_7584__bF_buf4), .C(_7303__bF_buf6_bF_buf3), .Y(_7805_) );
	OAI21X1 OAI21X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_7804_), .B(_7805_), .C(_7803_), .Y(_7806_) );
	NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf11), .B(_7806_), .Y(_7807_) );
	OAI21X1 OAI21X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf10), .B(_7799_), .C(_7807_), .Y(_6742__18_) );
	INVX1 INVX1_1334 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_19_), .Y(_7808_) );
	INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .Y(_7809_) );
	NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(biu_pc_18_), .C(_7789_), .Y(_7810_) );
	NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_7810_), .B(_7714_), .Y(_7811_) );
	XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_7811_), .B(_7809_), .Y(_7812_) );
	AOI21X1 AOI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(_7808_), .C(_7303__bF_buf5_bF_buf3), .Y(_7813_) );
	OAI21X1 OAI21X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7812_), .C(_7813_), .Y(_7814_) );
	NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf1), .B(_7586__bF_buf4), .Y(_7815_) );
	OAI21X1 OAI21X1_3414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_19_), .B(_7584__bF_buf3), .C(_7303__bF_buf4_bF_buf3), .Y(_7816_) );
	OAI21X1 OAI21X1_3415 ( .gnd(gnd), .vdd(vdd), .A(_7815_), .B(_7816_), .C(_7814_), .Y(_7817_) );
	NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf9), .B(_7817_), .Y(_7818_) );
	OAI21X1 OAI21X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf8), .B(_7808_), .C(_7818_), .Y(_6742__19_) );
	INVX1 INVX1_1335 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_20_), .Y(_7819_) );
	NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .B(_7811_), .Y(_7820_) );
	XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_7820_), .B(biu_pc_20_), .Y(_7821_) );
	AOI21X1 AOI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7819_), .C(_7303__bF_buf3_bF_buf3), .Y(_7822_) );
	OAI21X1 OAI21X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7821_), .C(_7822_), .Y(_7823_) );
	NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_7586__bF_buf3), .Y(_7824_) );
	OAI21X1 OAI21X1_3418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_20_), .B(_7584__bF_buf2), .C(_7303__bF_buf2), .Y(_7825_) );
	OAI21X1 OAI21X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_7824_), .B(_7825_), .C(_7823_), .Y(_7826_) );
	NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf7), .B(_7826_), .Y(_7827_) );
	OAI21X1 OAI21X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf6), .B(_7819_), .C(_7827_), .Y(_6742__20_) );
	INVX1 INVX1_1336 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_21_), .Y(_7828_) );
	NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .B(_7810_), .Y(_7829_) );
	NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_7829_), .C(_7725_), .Y(_7830_) );
	XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_7830_), .B(biu_pc_21_), .Y(_7831_) );
	AOI21X1 AOI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7828_), .C(_7303__bF_buf1), .Y(_7832_) );
	OAI21X1 OAI21X1_3421 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7831_), .C(_7832_), .Y(_7833_) );
	NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf1), .B(_7586__bF_buf2), .Y(_7834_) );
	OAI21X1 OAI21X1_3422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_21_), .B(_7584__bF_buf1), .C(_7303__bF_buf0), .Y(_7835_) );
	OAI21X1 OAI21X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_7834_), .B(_7835_), .C(_7833_), .Y(_7836_) );
	NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf5), .B(_7836_), .Y(_7837_) );
	OAI21X1 OAI21X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf4), .B(_7828_), .C(_7837_), .Y(_6742__21_) );
	INVX1 INVX1_1337 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_22_), .Y(_7838_) );
	INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .Y(_7839_) );
	INVX1 INVX1_1338 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .Y(_7840_) );
	NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_7840_), .B(_7830_), .Y(_7841_) );
	XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_7841_), .B(_7839_), .Y(_7842_) );
	AOI21X1 AOI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7838_), .C(_7303__bF_buf14_bF_buf2), .Y(_7843_) );
	OAI21X1 OAI21X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(_7842_), .C(_7843_), .Y(_7844_) );
	NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_7586__bF_buf1), .Y(_7845_) );
	OAI21X1 OAI21X1_3426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_22_), .B(_7584__bF_buf0), .C(_7303__bF_buf13_bF_buf2), .Y(_7846_) );
	OAI21X1 OAI21X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_7845_), .B(_7846_), .C(_7844_), .Y(_7847_) );
	NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf3), .B(_7847_), .Y(_7848_) );
	OAI21X1 OAI21X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf2), .B(_7838_), .C(_7848_), .Y(_6742__22_) );
	INVX1 INVX1_1339 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_23_), .Y(_7849_) );
	INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .Y(_7850_) );
	NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_7829_), .B(_7713_), .Y(_7851_) );
	NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(biu_pc_21_), .Y(_7852_) );
	INVX1 INVX1_1340 ( .gnd(gnd), .vdd(vdd), .A(_7852_), .Y(_7853_) );
	NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_7853_), .Y(_7854_) );
	OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_7630_), .B(_7854_), .Y(_7855_) );
	NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_7851_), .B(_7855_), .Y(_7856_) );
	XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_7856_), .B(_7850_), .Y(_7857_) );
	AOI21X1 AOI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7849_), .C(_7303__bF_buf12_bF_buf2), .Y(_7858_) );
	OAI21X1 OAI21X1_3429 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7857_), .C(_7858_), .Y(_7859_) );
	OAI21X1 OAI21X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf3), .B(_7309__bF_buf1), .C(csr_gpr_iu_csr_sepc_23_), .Y(_7860_) );
	OAI21X1 OAI21X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_7586__bF_buf0), .C(_7860_), .Y(_7861_) );
	AOI21X1 AOI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_7861_), .B(_7303__bF_buf11_bF_buf2), .C(rst_bF_buf40), .Y(_7862_) );
	AOI22X1 AOI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf39), .B(_7849_), .C(_7862_), .D(_7859_), .Y(_6742__23_) );
	INVX1 INVX1_1341 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_24_), .Y(_7863_) );
	NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .B(_7856_), .Y(_7864_) );
	XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_7864_), .B(biu_pc_24_), .Y(_7865_) );
	AOI21X1 AOI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7863_), .C(_7303__bF_buf10_bF_buf2), .Y(_7866_) );
	OAI21X1 OAI21X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7865_), .C(_7866_), .Y(_7867_) );
	NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_7586__bF_buf5), .Y(_7868_) );
	OAI21X1 OAI21X1_3433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_24_), .B(_7584__bF_buf5), .C(_7303__bF_buf9_bF_buf2), .Y(_7869_) );
	OAI21X1 OAI21X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_7868_), .B(_7869_), .C(_7867_), .Y(_7870_) );
	NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf1), .B(_7870_), .Y(_7871_) );
	OAI21X1 OAI21X1_3435 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf0), .B(_7863_), .C(_7871_), .Y(_6742__24_) );
	INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_25_), .Y(_7872_) );
	NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .B(biu_pc_24_), .Y(_7873_) );
	NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_7873_), .B(_7851_), .Y(_7874_) );
	INVX1 INVX1_1342 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .Y(_7875_) );
	NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_7875_), .B(_7854_), .Y(_7876_) );
	NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_7876_), .C(_7874_), .Y(_7877_) );
	INVX1 INVX1_1343 ( .gnd(gnd), .vdd(vdd), .A(_7854_), .Y(_7878_) );
	NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_7878_), .C(_7874_), .Y(_7879_) );
	NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_7875_), .B(_7879_), .Y(_7880_) );
	AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_7880_), .B(_7877_), .Y(_7881_) );
	AOI21X1 AOI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7872_), .C(_7303__bF_buf8_bF_buf2), .Y(_7882_) );
	OAI21X1 OAI21X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7881_), .C(_7882_), .Y(_7883_) );
	NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf1), .B(_7584__bF_buf4), .Y(_7884_) );
	OAI21X1 OAI21X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_7872_), .B(_7584__bF_buf3), .C(_7884_), .Y(_7885_) );
	AOI21X1 AOI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_7885_), .B(_7303__bF_buf7_bF_buf2), .C(rst_bF_buf38), .Y(_7886_) );
	AOI22X1 AOI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf37), .B(_7872_), .C(_7886_), .D(_7883_), .Y(_6742__25_) );
	OAI21X1 OAI21X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf2), .B(_7309__bF_buf0), .C(csr_gpr_iu_csr_sepc_26_), .Y(_7887_) );
	OAI21X1 OAI21X1_3439 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7586__bF_buf4), .C(_7887_), .Y(_7888_) );
	INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .Y(_7889_) );
	XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_7877_), .B(_7889_), .Y(_7890_) );
	AOI21X1 AOI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(csr_gpr_iu_csr_sepc_26_), .C(_7303__bF_buf6_bF_buf2), .Y(_7891_) );
	OAI21X1 OAI21X1_3440 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf6), .B(_7890_), .C(_7891_), .Y(_7892_) );
	OAI21X1 OAI21X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_7888_), .C(_7892_), .Y(_7893_) );
	NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf36), .B(csr_gpr_iu_csr_sepc_26_), .Y(_7894_) );
	OAI21X1 OAI21X1_3442 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf35), .B(_7893_), .C(_7894_), .Y(_6742__26_) );
	INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_27_), .Y(_7895_) );
	NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(_7877_), .Y(_7896_) );
	XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_7896_), .B(biu_pc_27_), .Y(_7897_) );
	NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_7897_), .Y(_7898_) );
	OAI21X1 OAI21X1_3443 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_27_), .B(_7428__bF_buf0), .C(_7898_), .Y(_7899_) );
	AOI21X1 AOI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_7586__bF_buf3), .B(_7895_), .C(_7304__bF_buf1), .Y(_7900_) );
	OAI21X1 OAI21X1_3444 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf1), .B(_7586__bF_buf2), .C(_7900_), .Y(_7901_) );
	OAI21X1 OAI21X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5_bF_buf2), .B(_7899_), .C(_7901_), .Y(_7902_) );
	NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf42), .B(_7902_), .Y(_7903_) );
	OAI21X1 OAI21X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf41), .B(_7895_), .C(_7903_), .Y(_6742__27_) );
	INVX1 INVX1_1344 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_28_), .Y(_7904_) );
	NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(biu_pc_27_), .Y(_7905_) );
	NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_7905_), .B(_7877_), .Y(_7906_) );
	XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_7906_), .B(biu_pc_28_), .Y(_7907_) );
	MUX2X1 MUX2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_7907_), .B(_7904_), .S(_7428__bF_buf8), .Y(_7908_) );
	OAI21X1 OAI21X1_3447 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf3), .C(_7908_), .Y(_7909_) );
	OAI21X1 OAI21X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf1), .B(_7309__bF_buf3), .C(csr_gpr_iu_csr_sepc_28_), .Y(_7910_) );
	OAI21X1 OAI21X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_7586__bF_buf1), .C(_7910_), .Y(_7911_) );
	AOI21X1 AOI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_7911_), .B(_7303__bF_buf4_bF_buf2), .C(rst_bF_buf34), .Y(_7912_) );
	AOI22X1 AOI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf33), .B(_7904_), .C(_7912_), .D(_7909_), .Y(_6742__28_) );
	INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_29_), .Y(_7913_) );
	NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(biu_pc_11_), .Y(_7914_) );
	NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7914_), .Y(_7915_) );
	NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .B(biu_pc_13_), .Y(_7916_) );
	NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_7916_), .B(_7775_), .Y(_7917_) );
	NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_7915_), .B(_7917_), .C(_7688_), .Y(_7918_) );
	NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .B(biu_pc_17_), .Y(_7919_) );
	NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(biu_pc_19_), .Y(_7920_) );
	NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_7919_), .B(_7920_), .Y(_7921_) );
	NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_7839_), .B(_7850_), .Y(_7922_) );
	NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_7853_), .B(_7922_), .C(_7921_), .Y(_7923_) );
	NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_7923_), .B(_7918_), .Y(_7924_) );
	NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .B(biu_pc_25_), .C(_7924_), .Y(_7925_) );
	NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_7905_), .B(_7925_), .Y(_7926_) );
	NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .B(_7620_), .C(_7926_), .Y(_7927_) );
	XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_7927_), .B(biu_pc_29_), .Y(_7928_) );
	AOI21X1 AOI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_7913_), .C(_7303__bF_buf3_bF_buf2), .Y(_7929_) );
	OAI21X1 OAI21X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf4), .B(_7928_), .C(_7929_), .Y(_7930_) );
	NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf1), .B(_7586__bF_buf0), .Y(_7931_) );
	OAI21X1 OAI21X1_3451 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_29_), .B(_7584__bF_buf2), .C(_7303__bF_buf2), .Y(_7932_) );
	OAI21X1 OAI21X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_7931_), .B(_7932_), .C(_7930_), .Y(_7933_) );
	NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf40), .B(_7933_), .Y(_7934_) );
	OAI21X1 OAI21X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf39), .B(_7913_), .C(_7934_), .Y(_6742__29_) );
	INVX1 INVX1_1345 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_30_), .Y(_7935_) );
	INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .Y(_7936_) );
	INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .Y(_7937_) );
	OAI21X1 OAI21X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_7936_), .B(_7927_), .C(_7937_), .Y(_7938_) );
	NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_7936_), .B(_7927_), .Y(_7939_) );
	NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(_7939_), .Y(_7940_) );
	AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_7940_), .B(_7938_), .Y(_7941_) );
	AOI21X1 AOI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf3), .B(_7935_), .C(_7303__bF_buf1), .Y(_7942_) );
	OAI21X1 OAI21X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf2), .B(_7941_), .C(_7942_), .Y(_7943_) );
	NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_7586__bF_buf5), .Y(_7944_) );
	OAI21X1 OAI21X1_3456 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_30_), .B(_7584__bF_buf1), .C(_7303__bF_buf0), .Y(_7945_) );
	OAI21X1 OAI21X1_3457 ( .gnd(gnd), .vdd(vdd), .A(_7944_), .B(_7945_), .C(_7943_), .Y(_7946_) );
	NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf38), .B(_7946_), .Y(_7947_) );
	OAI21X1 OAI21X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf37), .B(_7935_), .C(_7947_), .Y(_6742__30_) );
	INVX1 INVX1_1346 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_31_), .Y(_7948_) );
	XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_7940_), .B(biu_pc_31_), .Y(_7949_) );
	AOI21X1 AOI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf1), .B(_7948_), .C(_7303__bF_buf14_bF_buf1), .Y(_7950_) );
	OAI21X1 OAI21X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf0), .B(_7949_), .C(_7950_), .Y(_7951_) );
	OAI21X1 OAI21X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf0), .B(_7309__bF_buf2), .C(csr_gpr_iu_csr_sepc_31_), .Y(_7952_) );
	OAI21X1 OAI21X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_7278_), .B(_7586__bF_buf4), .C(_7952_), .Y(_7953_) );
	AOI21X1 AOI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_7953_), .B(_7303__bF_buf13_bF_buf1), .C(rst_bF_buf32), .Y(_7954_) );
	AOI22X1 AOI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf31), .B(_7948_), .C(_7954_), .D(_7951_), .Y(_6742__31_) );
	INVX1 INVX1_1347 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_0_), .Y(_7955_) );
	AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(csr_gpr_iu_csr_tval_0_), .Y(_7956_) );
	INVX1 INVX1_1348 ( .gnd(gnd), .vdd(vdd), .A(_7322_), .Y(_7957_) );
	NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_7431_), .Y(_7958_) );
	NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_7958_), .B(_7957_), .Y(_7959_) );
	INVX8 INVX8_65 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .Y(_7960_) );
	AOI22X1 AOI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_7956_), .C(_7325_), .D(_7960__bF_buf5), .Y(_7961_) );
	AOI21X1 AOI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .B(_7303__bF_buf12_bF_buf1), .C(_7438_), .Y(_7962_) );
	OAI22X1 OAI22X1_681 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_7962__bF_buf4), .C(rst_bF_buf30), .D(_7961_), .Y(_6751__0_) );
	INVX1 INVX1_1349 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_1_), .Y(_7963_) );
	AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf3), .B(csr_gpr_iu_csr_tval_1_), .Y(_7964_) );
	AOI22X1 AOI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7964_), .C(_7329_), .D(_7960__bF_buf4), .Y(_7965_) );
	OAI22X1 OAI22X1_682 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7962__bF_buf3), .C(rst_bF_buf29), .D(_7965_), .Y(_6751__1_) );
	INVX1 INVX1_1350 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_2_), .Y(_7966_) );
	AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf3), .B(csr_gpr_iu_csr_tval_2_), .Y(_7967_) );
	AOI22X1 AOI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7967_), .C(_7333_), .D(_7960__bF_buf3), .Y(_7968_) );
	OAI22X1 OAI22X1_683 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .B(_7962__bF_buf2), .C(rst_bF_buf28), .D(_7968_), .Y(_6751__2_) );
	INVX1 INVX1_1351 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_3_), .Y(_7969_) );
	AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf3), .B(csr_gpr_iu_csr_tval_3_), .Y(_7970_) );
	AOI22X1 AOI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7970_), .C(_7336_), .D(_7960__bF_buf2), .Y(_7971_) );
	OAI22X1 OAI22X1_684 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_7962__bF_buf1), .C(rst_bF_buf27), .D(_7971_), .Y(_6751__3_) );
	INVX1 INVX1_1352 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_4_), .Y(_7972_) );
	AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf3), .B(csr_gpr_iu_csr_tval_4_), .Y(_7973_) );
	AOI22X1 AOI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_7973_), .C(_7339_), .D(_7960__bF_buf1), .Y(_7974_) );
	OAI22X1 OAI22X1_685 ( .gnd(gnd), .vdd(vdd), .A(_7972_), .B(_7962__bF_buf0), .C(rst_bF_buf26), .D(_7974_), .Y(_6751__4_) );
	INVX1 INVX1_1353 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_5_), .Y(_7975_) );
	AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf3), .B(csr_gpr_iu_csr_tval_5_), .Y(_7976_) );
	AOI22X1 AOI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_7976_), .C(_7342_), .D(_7960__bF_buf0), .Y(_7977_) );
	OAI22X1 OAI22X1_686 ( .gnd(gnd), .vdd(vdd), .A(_7975_), .B(_7962__bF_buf4), .C(rst_bF_buf25), .D(_7977_), .Y(_6751__5_) );
	INVX1 INVX1_1354 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_6_), .Y(_7978_) );
	AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf3), .B(csr_gpr_iu_csr_tval_6_), .Y(_7979_) );
	AOI22X1 AOI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_7979_), .C(_7345_), .D(_7960__bF_buf5), .Y(_7980_) );
	OAI22X1 OAI22X1_687 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .B(_7962__bF_buf3), .C(rst_bF_buf24), .D(_7980_), .Y(_6751__6_) );
	INVX1 INVX1_1355 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_7_), .Y(_7981_) );
	AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf3), .B(csr_gpr_iu_csr_tval_7_), .Y(_7982_) );
	AOI22X1 AOI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_7982_), .C(_7348_), .D(_7960__bF_buf4), .Y(_7983_) );
	OAI22X1 OAI22X1_688 ( .gnd(gnd), .vdd(vdd), .A(_7981_), .B(_7962__bF_buf2), .C(rst_bF_buf23), .D(_7983_), .Y(_6751__7_) );
	INVX1 INVX1_1356 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_8_), .Y(_7984_) );
	AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf3), .B(csr_gpr_iu_csr_tval_8_), .Y(_7985_) );
	AOI22X1 AOI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_7985_), .C(_7351_), .D(_7960__bF_buf3), .Y(_7986_) );
	OAI22X1 OAI22X1_689 ( .gnd(gnd), .vdd(vdd), .A(_7984_), .B(_7962__bF_buf1), .C(rst_bF_buf22), .D(_7986_), .Y(_6751__8_) );
	INVX1 INVX1_1357 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_9_), .Y(_7987_) );
	AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf3), .B(csr_gpr_iu_csr_tval_9_), .Y(_7988_) );
	AOI22X1 AOI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_7988_), .C(_7354_), .D(_7960__bF_buf2), .Y(_7989_) );
	OAI22X1 OAI22X1_690 ( .gnd(gnd), .vdd(vdd), .A(_7987_), .B(_7962__bF_buf0), .C(rst_bF_buf21), .D(_7989_), .Y(_6751__9_) );
	INVX1 INVX1_1358 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_10_), .Y(_7990_) );
	AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(csr_gpr_iu_csr_tval_10_), .Y(_7991_) );
	AOI22X1 AOI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_7991_), .C(_7357_), .D(_7960__bF_buf1), .Y(_7992_) );
	OAI22X1 OAI22X1_691 ( .gnd(gnd), .vdd(vdd), .A(_7990_), .B(_7962__bF_buf4), .C(rst_bF_buf20), .D(_7992_), .Y(_6751__10_) );
	INVX1 INVX1_1359 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_11_), .Y(_7993_) );
	AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(csr_gpr_iu_csr_tval_11_), .Y(_7994_) );
	AOI22X1 AOI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_7994_), .C(_7360_), .D(_7960__bF_buf0), .Y(_7995_) );
	OAI22X1 OAI22X1_692 ( .gnd(gnd), .vdd(vdd), .A(_7993_), .B(_7962__bF_buf3), .C(rst_bF_buf19), .D(_7995_), .Y(_6751__11_) );
	INVX1 INVX1_1360 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_12_), .Y(_7996_) );
	AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(csr_gpr_iu_csr_tval_12_), .Y(_7997_) );
	AOI22X1 AOI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_7997_), .C(_7363_), .D(_7960__bF_buf5), .Y(_7998_) );
	OAI22X1 OAI22X1_693 ( .gnd(gnd), .vdd(vdd), .A(_7996_), .B(_7962__bF_buf2), .C(rst_bF_buf18), .D(_7998_), .Y(_6751__12_) );
	INVX1 INVX1_1361 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_13_), .Y(_7999_) );
	AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(csr_gpr_iu_csr_tval_13_), .Y(_8000_) );
	AOI22X1 AOI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_8000_), .C(_7492_), .D(_7960__bF_buf4), .Y(_8001_) );
	OAI22X1 OAI22X1_694 ( .gnd(gnd), .vdd(vdd), .A(_7999_), .B(_7962__bF_buf1), .C(rst_bF_buf17), .D(_8001_), .Y(_6751__13_) );
	INVX1 INVX1_1362 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_14_), .Y(_8002_) );
	AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(csr_gpr_iu_csr_tval_14_), .Y(_8003_) );
	AOI22X1 AOI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_8003_), .C(_7370_), .D(_7960__bF_buf3), .Y(_8004_) );
	OAI22X1 OAI22X1_695 ( .gnd(gnd), .vdd(vdd), .A(_8002_), .B(_7962__bF_buf0), .C(rst_bF_buf16), .D(_8004_), .Y(_6751__14_) );
	INVX1 INVX1_1363 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_15_), .Y(_8005_) );
	AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(csr_gpr_iu_csr_tval_15_), .Y(_8006_) );
	AOI22X1 AOI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_8006_), .C(_7501_), .D(_7960__bF_buf2), .Y(_8007_) );
	OAI22X1 OAI22X1_696 ( .gnd(gnd), .vdd(vdd), .A(_8005_), .B(_7962__bF_buf4), .C(rst_bF_buf15), .D(_8007_), .Y(_6751__15_) );
	INVX1 INVX1_1364 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_16_), .Y(_8008_) );
	AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf2), .B(csr_gpr_iu_csr_tval_16_), .Y(_8009_) );
	AOI22X1 AOI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_8009_), .C(_7376_), .D(_7960__bF_buf1), .Y(_8010_) );
	OAI22X1 OAI22X1_697 ( .gnd(gnd), .vdd(vdd), .A(_8008_), .B(_7962__bF_buf3), .C(rst_bF_buf14), .D(_8010_), .Y(_6751__16_) );
	INVX1 INVX1_1365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_17_), .Y(_8011_) );
	AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf2), .B(csr_gpr_iu_csr_tval_17_), .Y(_8012_) );
	AOI22X1 AOI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_8012_), .C(_7510_), .D(_7960__bF_buf0), .Y(_8013_) );
	OAI22X1 OAI22X1_698 ( .gnd(gnd), .vdd(vdd), .A(_8011_), .B(_7962__bF_buf2), .C(rst_bF_buf13), .D(_8013_), .Y(_6751__17_) );
	INVX1 INVX1_1366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_18_), .Y(_8014_) );
	AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf2), .B(csr_gpr_iu_csr_tval_18_), .Y(_8015_) );
	AOI22X1 AOI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_8015_), .C(_7382_), .D(_7960__bF_buf5), .Y(_8016_) );
	OAI22X1 OAI22X1_699 ( .gnd(gnd), .vdd(vdd), .A(_8014_), .B(_7962__bF_buf1), .C(rst_bF_buf12), .D(_8016_), .Y(_6751__18_) );
	INVX1 INVX1_1367 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_19_), .Y(_8017_) );
	AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf2), .B(csr_gpr_iu_csr_tval_19_), .Y(_8018_) );
	AOI22X1 AOI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_8018_), .C(_7519_), .D(_7960__bF_buf4), .Y(_8019_) );
	OAI22X1 OAI22X1_700 ( .gnd(gnd), .vdd(vdd), .A(_8017_), .B(_7962__bF_buf0), .C(rst_bF_buf11), .D(_8019_), .Y(_6751__19_) );
	INVX1 INVX1_1368 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_20_), .Y(_8020_) );
	AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf2), .B(csr_gpr_iu_csr_tval_20_), .Y(_8021_) );
	AOI22X1 AOI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_8021_), .C(_7388_), .D(_7960__bF_buf3), .Y(_8022_) );
	OAI22X1 OAI22X1_701 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_7962__bF_buf4), .C(rst_bF_buf10), .D(_8022_), .Y(_6751__20_) );
	INVX1 INVX1_1369 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_21_), .Y(_8023_) );
	AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf2), .B(csr_gpr_iu_csr_tval_21_), .Y(_8024_) );
	AOI22X1 AOI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_8024_), .C(_7528_), .D(_7960__bF_buf2), .Y(_8025_) );
	OAI22X1 OAI22X1_702 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_7962__bF_buf3), .C(rst_bF_buf9), .D(_8025_), .Y(_6751__21_) );
	INVX1 INVX1_1370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_22_), .Y(_8026_) );
	AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf2), .B(csr_gpr_iu_csr_tval_22_), .Y(_8027_) );
	AOI22X1 AOI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_8027_), .C(_7394_), .D(_7960__bF_buf1), .Y(_8028_) );
	OAI22X1 OAI22X1_703 ( .gnd(gnd), .vdd(vdd), .A(_8026_), .B(_7962__bF_buf2), .C(rst_bF_buf8), .D(_8028_), .Y(_6751__22_) );
	INVX1 INVX1_1371 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_23_), .Y(_8029_) );
	AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf2), .B(csr_gpr_iu_csr_tval_23_), .Y(_8030_) );
	AOI22X1 AOI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf2), .B(_8030_), .C(_7537_), .D(_7960__bF_buf0), .Y(_8031_) );
	OAI22X1 OAI22X1_704 ( .gnd(gnd), .vdd(vdd), .A(_8029_), .B(_7962__bF_buf1), .C(rst_bF_buf7), .D(_8031_), .Y(_6751__23_) );
	INVX1 INVX1_1372 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_24_), .Y(_8032_) );
	AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf2), .B(csr_gpr_iu_csr_tval_24_), .Y(_8033_) );
	AOI22X1 AOI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf1), .B(_8033_), .C(_7400_), .D(_7960__bF_buf5), .Y(_8034_) );
	OAI22X1 OAI22X1_705 ( .gnd(gnd), .vdd(vdd), .A(_8032_), .B(_7962__bF_buf0), .C(rst_bF_buf6), .D(_8034_), .Y(_6751__24_) );
	INVX1 INVX1_1373 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_25_), .Y(_8035_) );
	AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(csr_gpr_iu_csr_tval_25_), .Y(_8036_) );
	AOI22X1 AOI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf0), .B(_8036_), .C(_7546_), .D(_7960__bF_buf4), .Y(_8037_) );
	OAI22X1 OAI22X1_706 ( .gnd(gnd), .vdd(vdd), .A(_8035_), .B(_7962__bF_buf4), .C(rst_bF_buf5), .D(_8037_), .Y(_6751__25_) );
	INVX1 INVX1_1374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_26_), .Y(_8038_) );
	AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(csr_gpr_iu_csr_tval_26_), .Y(_8039_) );
	AOI22X1 AOI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_8039_), .C(_7406_), .D(_7960__bF_buf3), .Y(_8040_) );
	OAI22X1 OAI22X1_707 ( .gnd(gnd), .vdd(vdd), .A(_8038_), .B(_7962__bF_buf3), .C(rst_bF_buf4), .D(_8040_), .Y(_6751__26_) );
	INVX1 INVX1_1375 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_27_), .Y(_8041_) );
	AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(csr_gpr_iu_csr_tval_27_), .Y(_8042_) );
	AOI22X1 AOI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf7), .B(_8042_), .C(_7556_), .D(_7960__bF_buf2), .Y(_8043_) );
	OAI22X1 OAI22X1_708 ( .gnd(gnd), .vdd(vdd), .A(_8041_), .B(_7962__bF_buf2), .C(rst_bF_buf3), .D(_8043_), .Y(_6751__27_) );
	INVX1 INVX1_1376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_28_), .Y(_8044_) );
	AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(csr_gpr_iu_csr_tval_28_), .Y(_8045_) );
	AOI22X1 AOI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf6), .B(_8045_), .C(_7412_), .D(_7960__bF_buf1), .Y(_8046_) );
	OAI22X1 OAI22X1_709 ( .gnd(gnd), .vdd(vdd), .A(_8044_), .B(_7962__bF_buf1), .C(rst_bF_buf2), .D(_8046_), .Y(_6751__28_) );
	INVX1 INVX1_1377 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_29_), .Y(_8047_) );
	AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(csr_gpr_iu_csr_tval_29_), .Y(_8048_) );
	AOI22X1 AOI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf5), .B(_8048_), .C(_7565_), .D(_7960__bF_buf0), .Y(_8049_) );
	OAI22X1 OAI22X1_710 ( .gnd(gnd), .vdd(vdd), .A(_8047_), .B(_7962__bF_buf0), .C(rst_bF_buf1), .D(_8049_), .Y(_6751__29_) );
	INVX1 INVX1_1378 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_30_), .Y(_8050_) );
	AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(csr_gpr_iu_csr_tval_30_), .Y(_8051_) );
	AOI22X1 AOI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf4), .B(_8051_), .C(_7417_), .D(_7960__bF_buf5), .Y(_8052_) );
	OAI22X1 OAI22X1_711 ( .gnd(gnd), .vdd(vdd), .A(_8050_), .B(_7962__bF_buf4), .C(rst_bF_buf0), .D(_8052_), .Y(_6751__30_) );
	INVX1 INVX1_1379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_31_), .Y(_8053_) );
	AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf1), .B(csr_gpr_iu_csr_tval_31_), .Y(_8054_) );
	AOI22X1 AOI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf3), .B(_8054_), .C(_7574_), .D(_7960__bF_buf4), .Y(_8055_) );
	OAI22X1 OAI22X1_712 ( .gnd(gnd), .vdd(vdd), .A(_8053_), .B(_7962__bF_buf3), .C(rst_bF_buf70), .D(_8055_), .Y(_6751__31_) );
	NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf2), .B(biu_ins_27_bF_buf3), .Y(_8056_) );
	NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_8056_), .Y(_8057_) );
	NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .B(_6779_), .Y(_8058_) );
	NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_7580_), .B(_8058_), .Y(_8059_) );
	NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_8057_), .B(_8059_), .Y(_8060_) );
	NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_8060_), .B(_7308_), .Y(_8061_) );
	INVX8 INVX8_66 ( .gnd(gnd), .vdd(vdd), .A(_8061_), .Y(_8062_) );
	NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11_bF_buf1), .B(_8062__bF_buf5), .Y(_8063_) );
	AOI22X1 AOI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8062__bF_buf4), .C(csr_gpr_iu_csr_stvec_0_), .D(_8063__bF_buf5), .Y(_8064_) );
	NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf69), .B(_8064_), .Y(_6752__0_) );
	AOI22X1 AOI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8062__bF_buf3), .C(csr_gpr_iu_csr_stvec_1_), .D(_8063__bF_buf4), .Y(_8065_) );
	NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_8065_), .Y(_6752__1_) );
	AOI22X1 AOI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8062__bF_buf2), .C(csr_gpr_iu_csr_stvec_2_), .D(_8063__bF_buf3), .Y(_8066_) );
	NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf67), .B(_8066_), .Y(_6752__2_) );
	AOI22X1 AOI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8062__bF_buf1), .C(csr_gpr_iu_csr_stvec_3_), .D(_8063__bF_buf2), .Y(_8067_) );
	NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf66), .B(_8067_), .Y(_6752__3_) );
	AOI22X1 AOI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8062__bF_buf0), .C(csr_gpr_iu_csr_stvec_4_), .D(_8063__bF_buf1), .Y(_8068_) );
	NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf65), .B(_8068_), .Y(_6752__4_) );
	AOI22X1 AOI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8062__bF_buf5), .C(csr_gpr_iu_csr_stvec_5_), .D(_8063__bF_buf0), .Y(_8069_) );
	NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf64), .B(_8069_), .Y(_6752__5_) );
	AOI22X1 AOI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8062__bF_buf4), .C(csr_gpr_iu_csr_stvec_6_), .D(_8063__bF_buf5), .Y(_8070_) );
	NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf63), .B(_8070_), .Y(_6752__6_) );
	AOI22X1 AOI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8062__bF_buf3), .C(csr_gpr_iu_csr_stvec_7_), .D(_8063__bF_buf4), .Y(_8071_) );
	NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf62), .B(_8071_), .Y(_6752__7_) );
	AOI22X1 AOI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8062__bF_buf2), .C(csr_gpr_iu_csr_stvec_8_), .D(_8063__bF_buf3), .Y(_8072_) );
	NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf61), .B(_8072_), .Y(_6752__8_) );
	AOI22X1 AOI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8062__bF_buf1), .C(csr_gpr_iu_csr_stvec_9_), .D(_8063__bF_buf2), .Y(_8073_) );
	NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf60), .B(_8073_), .Y(_6752__9_) );
	AOI22X1 AOI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8062__bF_buf0), .C(csr_gpr_iu_csr_stvec_10_), .D(_8063__bF_buf1), .Y(_8074_) );
	NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf59), .B(_8074_), .Y(_6752__10_) );
	AOI22X1 AOI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8062__bF_buf5), .C(csr_gpr_iu_csr_stvec_11_), .D(_8063__bF_buf0), .Y(_8075_) );
	NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf58), .B(_8075_), .Y(_6752__11_) );
	AOI22X1 AOI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8062__bF_buf4), .C(csr_gpr_iu_csr_stvec_12_), .D(_8063__bF_buf5), .Y(_8076_) );
	NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf57), .B(_8076_), .Y(_6752__12_) );
	INVX1 INVX1_1380 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_13_), .Y(_8077_) );
	OAI21X1 OAI21X1_3462 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf1), .B(_8063__bF_buf4), .C(_6879__bF_buf36), .Y(_8078_) );
	AOI21X1 AOI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .B(_8063__bF_buf3), .C(_8078_), .Y(_6752__13_) );
	AOI22X1 AOI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf2), .B(csr_gpr_iu_csr_stvec_14_), .C(_7370_), .D(_8062__bF_buf3), .Y(_8079_) );
	NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf56), .B(_8079_), .Y(_6752__14_) );
	INVX1 INVX1_1381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_15_), .Y(_8080_) );
	OAI21X1 OAI21X1_3463 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf2), .B(_8063__bF_buf1), .C(_6879__bF_buf35), .Y(_8081_) );
	AOI21X1 AOI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_8063__bF_buf0), .C(_8081_), .Y(_6752__15_) );
	AOI22X1 AOI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf5), .B(csr_gpr_iu_csr_stvec_16_), .C(_7376_), .D(_8062__bF_buf2), .Y(_8082_) );
	NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf55), .B(_8082_), .Y(_6752__16_) );
	INVX1 INVX1_1382 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_17_), .Y(_8083_) );
	OAI21X1 OAI21X1_3464 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf3), .B(_8063__bF_buf4), .C(_6879__bF_buf34), .Y(_8084_) );
	AOI21X1 AOI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_8063__bF_buf3), .C(_8084_), .Y(_6752__17_) );
	AOI22X1 AOI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf2), .B(csr_gpr_iu_csr_stvec_18_), .C(_7382_), .D(_8062__bF_buf1), .Y(_8085_) );
	NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf54), .B(_8085_), .Y(_6752__18_) );
	INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_19_), .Y(_8086_) );
	OAI21X1 OAI21X1_3465 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf0), .B(_8063__bF_buf1), .C(_6879__bF_buf33), .Y(_8087_) );
	AOI21X1 AOI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_8086_), .B(_8063__bF_buf0), .C(_8087_), .Y(_6752__19_) );
	AOI22X1 AOI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf5), .B(csr_gpr_iu_csr_stvec_20_), .C(_7388_), .D(_8062__bF_buf0), .Y(_8088_) );
	NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf53), .B(_8088_), .Y(_6752__20_) );
	INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_21_), .Y(_8089_) );
	OAI21X1 OAI21X1_3466 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf0), .B(_8063__bF_buf4), .C(_6879__bF_buf32), .Y(_8090_) );
	AOI21X1 AOI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .B(_8063__bF_buf3), .C(_8090_), .Y(_6752__21_) );
	AOI22X1 AOI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf2), .B(csr_gpr_iu_csr_stvec_22_), .C(_7394_), .D(_8062__bF_buf5), .Y(_8091_) );
	NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf52), .B(_8091_), .Y(_6752__22_) );
	INVX1 INVX1_1383 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_23_), .Y(_8092_) );
	OAI21X1 OAI21X1_3467 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf2), .B(_8063__bF_buf1), .C(_6879__bF_buf31), .Y(_8093_) );
	AOI21X1 AOI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_8063__bF_buf0), .C(_8093_), .Y(_6752__23_) );
	AOI22X1 AOI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf5), .B(csr_gpr_iu_csr_stvec_24_), .C(_7400_), .D(_8062__bF_buf4), .Y(_8094_) );
	NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf51), .B(_8094_), .Y(_6752__24_) );
	INVX1 INVX1_1384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_25_), .Y(_8095_) );
	OAI21X1 OAI21X1_3468 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf0), .B(_8063__bF_buf4), .C(_6879__bF_buf30), .Y(_8096_) );
	AOI21X1 AOI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_8095_), .B(_8063__bF_buf3), .C(_8096_), .Y(_6752__25_) );
	AOI22X1 AOI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf2), .B(csr_gpr_iu_csr_stvec_26_), .C(_7406_), .D(_8062__bF_buf3), .Y(_8097_) );
	NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf50), .B(_8097_), .Y(_6752__26_) );
	INVX1 INVX1_1385 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_27_), .Y(_8098_) );
	OAI21X1 OAI21X1_3469 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf0), .B(_8063__bF_buf1), .C(_6879__bF_buf29), .Y(_8099_) );
	AOI21X1 AOI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_8063__bF_buf0), .C(_8099_), .Y(_6752__27_) );
	AOI22X1 AOI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf5), .B(csr_gpr_iu_csr_stvec_28_), .C(_7412_), .D(_8062__bF_buf2), .Y(_8100_) );
	NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf49), .B(_8100_), .Y(_6752__28_) );
	INVX1 INVX1_1386 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_29_), .Y(_8101_) );
	OAI21X1 OAI21X1_3470 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf0), .B(_8063__bF_buf4), .C(_6879__bF_buf28), .Y(_8102_) );
	AOI21X1 AOI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_8101_), .B(_8063__bF_buf3), .C(_8102_), .Y(_6752__29_) );
	AOI22X1 AOI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(_8063__bF_buf2), .B(csr_gpr_iu_csr_stvec_30_), .C(_7417_), .D(_8062__bF_buf1), .Y(_8103_) );
	NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf48), .B(_8103_), .Y(_6752__30_) );
	INVX1 INVX1_1387 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_31_), .Y(_8104_) );
	OAI21X1 OAI21X1_3471 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf2), .B(_8063__bF_buf1), .C(_6879__bF_buf27), .Y(_8105_) );
	AOI21X1 AOI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_8104_), .B(_8063__bF_buf0), .C(_8105_), .Y(_6752__31_) );
	INVX1 INVX1_1388 ( .gnd(gnd), .vdd(vdd), .A(_7958_), .Y(_8106_) );
	INVX1 INVX1_1389 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf2), .Y(_8107_) );
	NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_8107_), .Y(_8108_) );
	INVX1 INVX1_1390 ( .gnd(gnd), .vdd(vdd), .A(_8108_), .Y(_8109_) );
	NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_7305_), .B(_8109_), .Y(_8110_) );
	INVX8 INVX8_67 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .Y(_8111_) );
	NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_8106_), .B(_8111__bF_buf5), .Y(_8112_) );
	NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf1), .B(_6799_), .Y(_8113_) );
	AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .B(biu_ins_25_bF_buf3), .Y(_8114_) );
	AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_8113_), .B(_8114_), .Y(_8115_) );
	NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_8112_), .Y(_8116_) );
	INVX8 INVX8_68 ( .gnd(gnd), .vdd(vdd), .A(_8116_), .Y(_8117_) );
	NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf1), .B(_8117__bF_buf6), .Y(_8118_) );
	AOI22X1 AOI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8117__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr3_0_), .D(_8118__bF_buf5), .Y(_8119_) );
	NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf47), .B(_8119_), .Y(_6737__0_) );
	AOI22X1 AOI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8117__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr3_1_), .D(_8118__bF_buf4), .Y(_8120_) );
	NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf46), .B(_8120_), .Y(_6737__1_) );
	AOI22X1 AOI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8117__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_2_), .D(_8118__bF_buf3), .Y(_8121_) );
	NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf45), .B(_8121_), .Y(_6737__2_) );
	AOI22X1 AOI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr3_3_), .D(_8118__bF_buf2), .Y(_8122_) );
	NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf44), .B(_8122_), .Y(_6737__3_) );
	AOI22X1 AOI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8117__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_4_), .D(_8118__bF_buf1), .Y(_8123_) );
	NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf43), .B(_8123_), .Y(_6737__4_) );
	AOI22X1 AOI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8117__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr3_5_), .D(_8118__bF_buf0), .Y(_8124_) );
	NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf42), .B(_8124_), .Y(_6737__5_) );
	AOI22X1 AOI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8117__bF_buf6), .C(csr_gpr_iu_csr_pmpaddr3_6_), .D(_8118__bF_buf5), .Y(_8125_) );
	NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf41), .B(_8125_), .Y(_6737__6_) );
	AOI22X1 AOI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8117__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr3_7_), .D(_8118__bF_buf4), .Y(_8126_) );
	NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf40), .B(_8126_), .Y(_6737__7_) );
	AOI22X1 AOI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8117__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr3_8_), .D(_8118__bF_buf3), .Y(_8127_) );
	NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf39), .B(_8127_), .Y(_6737__8_) );
	AOI22X1 AOI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8117__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_9_), .D(_8118__bF_buf2), .Y(_8128_) );
	NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf38), .B(_8128_), .Y(_6737__9_) );
	AOI22X1 AOI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr3_10_), .D(_8118__bF_buf1), .Y(_8129_) );
	NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf37), .B(_8129_), .Y(_6737__10_) );
	AOI22X1 AOI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8117__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_11_), .D(_8118__bF_buf0), .Y(_8130_) );
	NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf36), .B(_8130_), .Y(_6737__11_) );
	AOI22X1 AOI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8117__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr3_12_), .D(_8118__bF_buf5), .Y(_8131_) );
	NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf35), .B(_8131_), .Y(_6737__12_) );
	INVX1 INVX1_1391 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_13_), .Y(_8132_) );
	OAI21X1 OAI21X1_3472 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf0), .B(_8118__bF_buf4), .C(_6879__bF_buf26), .Y(_8133_) );
	AOI21X1 AOI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_8132_), .B(_8118__bF_buf3), .C(_8133_), .Y(_6737__13_) );
	AOI22X1 AOI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8117__bF_buf6), .C(csr_gpr_iu_csr_pmpaddr3_14_), .D(_8118__bF_buf2), .Y(_8134_) );
	NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf34), .B(_8134_), .Y(_6737__14_) );
	INVX1 INVX1_1392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_15_), .Y(_8135_) );
	OAI21X1 OAI21X1_3473 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf1), .B(_8118__bF_buf1), .C(_6879__bF_buf25), .Y(_8136_) );
	AOI21X1 AOI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_8135_), .B(_8118__bF_buf0), .C(_8136_), .Y(_6737__15_) );
	AOI22X1 AOI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_8117__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr3_16_), .D(_8118__bF_buf5), .Y(_8137_) );
	NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf33), .B(_8137_), .Y(_6737__16_) );
	INVX1 INVX1_1393 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_17_), .Y(_8138_) );
	OAI21X1 OAI21X1_3474 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf2), .B(_8118__bF_buf4), .C(_6879__bF_buf24), .Y(_8139_) );
	AOI21X1 AOI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_8138_), .B(_8118__bF_buf3), .C(_8139_), .Y(_6737__17_) );
	AOI22X1 AOI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8117__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr3_18_), .D(_8118__bF_buf2), .Y(_8140_) );
	NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf32), .B(_8140_), .Y(_6737__18_) );
	INVX1 INVX1_1394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_19_), .Y(_8141_) );
	OAI21X1 OAI21X1_3475 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_8118__bF_buf1), .C(_6879__bF_buf23), .Y(_8142_) );
	AOI21X1 AOI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .B(_8118__bF_buf0), .C(_8142_), .Y(_6737__19_) );
	AOI22X1 AOI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8117__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_20_), .D(_8118__bF_buf5), .Y(_8143_) );
	NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf31), .B(_8143_), .Y(_6737__20_) );
	INVX1 INVX1_1395 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_21_), .Y(_8144_) );
	OAI21X1 OAI21X1_3476 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_8118__bF_buf4), .C(_6879__bF_buf22), .Y(_8145_) );
	AOI21X1 AOI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_8144_), .B(_8118__bF_buf3), .C(_8145_), .Y(_6737__21_) );
	AOI22X1 AOI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr3_22_), .D(_8118__bF_buf2), .Y(_8146_) );
	NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf30), .B(_8146_), .Y(_6737__22_) );
	INVX1 INVX1_1396 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_23_), .Y(_8147_) );
	OAI21X1 OAI21X1_3477 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf1), .B(_8118__bF_buf1), .C(_6879__bF_buf21), .Y(_8148_) );
	AOI21X1 AOI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_8147_), .B(_8118__bF_buf0), .C(_8148_), .Y(_6737__23_) );
	AOI22X1 AOI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_8117__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_24_), .D(_8118__bF_buf5), .Y(_8149_) );
	NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf29), .B(_8149_), .Y(_6737__24_) );
	INVX1 INVX1_1397 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_25_), .Y(_8150_) );
	OAI21X1 OAI21X1_3478 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_8118__bF_buf4), .C(_6879__bF_buf20), .Y(_8151_) );
	AOI21X1 AOI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_8150_), .B(_8118__bF_buf3), .C(_8151_), .Y(_6737__25_) );
	AOI22X1 AOI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(_7406_), .B(_8117__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr3_26_), .D(_8118__bF_buf2), .Y(_8152_) );
	NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf28), .B(_8152_), .Y(_6737__26_) );
	INVX1 INVX1_1398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_27_), .Y(_8153_) );
	OAI21X1 OAI21X1_3479 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_8118__bF_buf1), .C(_6879__bF_buf19), .Y(_8154_) );
	AOI21X1 AOI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .B(_8118__bF_buf0), .C(_8154_), .Y(_6737__27_) );
	AOI22X1 AOI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8117__bF_buf6), .C(csr_gpr_iu_csr_pmpaddr3_28_), .D(_8118__bF_buf5), .Y(_8155_) );
	NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf27), .B(_8155_), .Y(_6737__28_) );
	INVX1 INVX1_1399 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_29_), .Y(_8156_) );
	OAI21X1 OAI21X1_3480 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_8118__bF_buf4), .C(_6879__bF_buf18), .Y(_8157_) );
	AOI21X1 AOI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_8156_), .B(_8118__bF_buf3), .C(_8157_), .Y(_6737__29_) );
	AOI22X1 AOI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8117__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr3_30_), .D(_8118__bF_buf2), .Y(_8158_) );
	NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf26), .B(_8158_), .Y(_6737__30_) );
	INVX1 INVX1_1400 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_31_), .Y(_8159_) );
	OAI21X1 OAI21X1_3481 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf1), .B(_8118__bF_buf1), .C(_6879__bF_buf17), .Y(_8160_) );
	AOI21X1 AOI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_8159_), .B(_8118__bF_buf0), .C(_8160_), .Y(_6737__31_) );
	NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_7432_), .B(_8111__bF_buf4), .Y(_8161_) );
	NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_8161_), .Y(_8162_) );
	OAI21X1 OAI21X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf1), .B(_8162__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_0_), .Y(_8163_) );
	NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_7433_), .Y(_8164_) );
	NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_8164_), .Y(_8165_) );
	NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf4), .B(_7325_), .Y(_8166_) );
	AOI21X1 AOI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_8163_), .B(_8166_), .C(rst_bF_buf25), .Y(_6736__0_) );
	OAI21X1 OAI21X1_3483 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf1), .B(_8162__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_1_), .Y(_8167_) );
	NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf3), .B(_7329_), .Y(_8168_) );
	AOI21X1 AOI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_8167_), .B(_8168_), .C(rst_bF_buf24), .Y(_6736__1_) );
	OAI21X1 OAI21X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf1), .B(_8162__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr2_2_), .Y(_8169_) );
	NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(_7333_), .Y(_8170_) );
	AOI21X1 AOI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_8169_), .B(_8170_), .C(rst_bF_buf23), .Y(_6736__2_) );
	OAI21X1 OAI21X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf1), .B(_8162__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr2_3_), .Y(_8171_) );
	NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf1), .B(_7336_), .Y(_8172_) );
	AOI21X1 AOI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(_8172_), .C(rst_bF_buf22), .Y(_6736__3_) );
	OAI21X1 OAI21X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf1), .B(_8162__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr2_4_), .Y(_8173_) );
	NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf0), .B(_7339_), .Y(_8174_) );
	AOI21X1 AOI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_8173_), .B(_8174_), .C(rst_bF_buf21), .Y(_6736__4_) );
	OAI21X1 OAI21X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf1), .B(_8162__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_5_), .Y(_8175_) );
	NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf4), .B(_7342_), .Y(_8176_) );
	AOI21X1 AOI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_8175_), .B(_8176_), .C(rst_bF_buf20), .Y(_6736__5_) );
	OAI21X1 OAI21X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf1), .B(_8162__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_6_), .Y(_8177_) );
	NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf3), .B(_7345_), .Y(_8178_) );
	AOI21X1 AOI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_8177_), .B(_8178_), .C(rst_bF_buf19), .Y(_6736__6_) );
	OAI21X1 OAI21X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf1), .B(_8162__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr2_7_), .Y(_8179_) );
	NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(_7348_), .Y(_8180_) );
	AOI21X1 AOI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_8179_), .B(_8180_), .C(rst_bF_buf18), .Y(_6736__7_) );
	OAI21X1 OAI21X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_8162__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr2_8_), .Y(_8181_) );
	NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf1), .B(_7351_), .Y(_8182_) );
	AOI21X1 AOI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_8181_), .B(_8182_), .C(rst_bF_buf17), .Y(_6736__8_) );
	OAI21X1 OAI21X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_8162__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr2_9_), .Y(_8183_) );
	NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf0), .B(_7354_), .Y(_8184_) );
	AOI21X1 AOI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_8183_), .B(_8184_), .C(rst_bF_buf16), .Y(_6736__9_) );
	OAI21X1 OAI21X1_3492 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_8162__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_10_), .Y(_8185_) );
	NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf4), .B(_7357_), .Y(_8186_) );
	AOI21X1 AOI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_8185_), .B(_8186_), .C(rst_bF_buf15), .Y(_6736__10_) );
	OAI21X1 OAI21X1_3493 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_8162__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_11_), .Y(_8187_) );
	NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf3), .B(_7360_), .Y(_8188_) );
	AOI21X1 AOI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_8187_), .B(_8188_), .C(rst_bF_buf14), .Y(_6736__11_) );
	OAI21X1 OAI21X1_3494 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_8162__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr2_12_), .Y(_8189_) );
	NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(_7363_), .Y(_8190_) );
	AOI21X1 AOI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_8189_), .B(_8190_), .C(rst_bF_buf13), .Y(_6736__12_) );
	INVX1 INVX1_1401 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_13_), .Y(_8191_) );
	NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9_bF_buf1), .B(_8165__bF_buf1), .Y(_8192_) );
	OAI21X1 OAI21X1_3495 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_8192__bF_buf3), .C(_6879__bF_buf16), .Y(_8193_) );
	AOI21X1 AOI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_8192__bF_buf2), .C(_8193_), .Y(_6736__13_) );
	OAI21X1 OAI21X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(_8162__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr2_14_), .Y(_8194_) );
	NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf0), .B(_7370_), .Y(_8195_) );
	AOI21X1 AOI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_8194_), .B(_8195_), .C(rst_bF_buf12), .Y(_6736__14_) );
	INVX1 INVX1_1402 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_15_), .Y(_8196_) );
	OAI21X1 OAI21X1_3497 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf0), .B(_8192__bF_buf1), .C(_6879__bF_buf15), .Y(_8197_) );
	AOI21X1 AOI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_8196_), .B(_8192__bF_buf0), .C(_8197_), .Y(_6736__15_) );
	OAI21X1 OAI21X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf0), .B(_8162__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr2_16_), .Y(_8198_) );
	NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf4), .B(_7376_), .Y(_8199_) );
	AOI21X1 AOI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_8198_), .B(_8199_), .C(rst_bF_buf11), .Y(_6736__16_) );
	INVX1 INVX1_1403 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_17_), .Y(_8200_) );
	OAI21X1 OAI21X1_3499 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf1), .B(_8192__bF_buf3), .C(_6879__bF_buf14), .Y(_8201_) );
	AOI21X1 AOI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_8200_), .B(_8192__bF_buf2), .C(_8201_), .Y(_6736__17_) );
	OAI21X1 OAI21X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf0), .B(_8162__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_18_), .Y(_8202_) );
	NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf3), .B(_7382_), .Y(_8203_) );
	AOI21X1 AOI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_8202_), .B(_8203_), .C(rst_bF_buf10), .Y(_6736__18_) );
	INVX1 INVX1_1404 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_19_), .Y(_8204_) );
	OAI21X1 OAI21X1_3501 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf2), .B(_8192__bF_buf1), .C(_6879__bF_buf13), .Y(_8205_) );
	AOI21X1 AOI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_8204_), .B(_8192__bF_buf0), .C(_8205_), .Y(_6736__19_) );
	OAI21X1 OAI21X1_3502 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf0), .B(_8162__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_20_), .Y(_8206_) );
	NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(_7388_), .Y(_8207_) );
	AOI21X1 AOI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_8206_), .B(_8207_), .C(rst_bF_buf9), .Y(_6736__20_) );
	INVX1 INVX1_1405 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_21_), .Y(_8208_) );
	OAI21X1 OAI21X1_3503 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf2), .B(_8192__bF_buf3), .C(_6879__bF_buf12), .Y(_8209_) );
	AOI21X1 AOI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_8208_), .B(_8192__bF_buf2), .C(_8209_), .Y(_6736__21_) );
	OAI21X1 OAI21X1_3504 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf0), .B(_8162__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr2_22_), .Y(_8210_) );
	NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf1), .B(_7394_), .Y(_8211_) );
	AOI21X1 AOI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_8210_), .B(_8211_), .C(rst_bF_buf8), .Y(_6736__22_) );
	INVX1 INVX1_1406 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_23_), .Y(_8212_) );
	OAI21X1 OAI21X1_3505 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf0), .B(_8192__bF_buf1), .C(_6879__bF_buf11), .Y(_8213_) );
	AOI21X1 AOI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8192__bF_buf0), .C(_8213_), .Y(_6736__23_) );
	OAI21X1 OAI21X1_3506 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf0), .B(_8162__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr2_24_), .Y(_8214_) );
	NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf0), .B(_7400_), .Y(_8215_) );
	AOI21X1 AOI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_8214_), .B(_8215_), .C(rst_bF_buf7), .Y(_6736__24_) );
	INVX1 INVX1_1407 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_25_), .Y(_8216_) );
	OAI21X1 OAI21X1_3507 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf2), .B(_8192__bF_buf3), .C(_6879__bF_buf10), .Y(_8217_) );
	AOI21X1 AOI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_8216_), .B(_8192__bF_buf2), .C(_8217_), .Y(_6736__25_) );
	OAI21X1 OAI21X1_3508 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf0), .B(_8162__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr2_26_), .Y(_8218_) );
	NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf4), .B(_7406_), .Y(_8219_) );
	AOI21X1 AOI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_8218_), .B(_8219_), .C(rst_bF_buf6), .Y(_6736__26_) );
	INVX1 INVX1_1408 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_27_), .Y(_8220_) );
	OAI21X1 OAI21X1_3509 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf2), .B(_8192__bF_buf1), .C(_6879__bF_buf9), .Y(_8221_) );
	AOI21X1 AOI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_8220_), .B(_8192__bF_buf0), .C(_8221_), .Y(_6736__27_) );
	OAI21X1 OAI21X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf0), .B(_8162__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_28_), .Y(_8222_) );
	NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf3), .B(_7412_), .Y(_8223_) );
	AOI21X1 AOI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_8222_), .B(_8223_), .C(rst_bF_buf5), .Y(_6736__28_) );
	INVX1 INVX1_1409 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_29_), .Y(_8224_) );
	OAI21X1 OAI21X1_3511 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf2), .B(_8192__bF_buf3), .C(_6879__bF_buf8), .Y(_8225_) );
	AOI21X1 AOI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_8224_), .B(_8192__bF_buf2), .C(_8225_), .Y(_6736__29_) );
	OAI21X1 OAI21X1_3512 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf0), .B(_8162__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_30_), .Y(_8226_) );
	NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(_7417_), .Y(_8227_) );
	AOI21X1 AOI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_8226_), .B(_8227_), .C(rst_bF_buf4), .Y(_6736__30_) );
	INVX1 INVX1_1410 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_31_), .Y(_8228_) );
	OAI21X1 OAI21X1_3513 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf0), .B(_8192__bF_buf1), .C(_6879__bF_buf7), .Y(_8229_) );
	AOI21X1 AOI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_8228_), .B(_8192__bF_buf0), .C(_8229_), .Y(_6736__31_) );
	NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_7582_), .B(_8110_), .Y(_8230_) );
	INVX1 INVX1_1411 ( .gnd(gnd), .vdd(vdd), .A(_8230_), .Y(_8231_) );
	NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_8231_), .Y(_8232_) );
	INVX8 INVX8_69 ( .gnd(gnd), .vdd(vdd), .A(_8232_), .Y(_8233_) );
	NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf0), .B(_8232_), .Y(_8234_) );
	INVX8 INVX8_70 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .Y(_8235_) );
	AOI22X1 AOI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8233__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr1_0_), .D(_8235__bF_buf5), .Y(_8236_) );
	NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_8236_), .Y(_6735__0_) );
	AOI22X1 AOI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr1_1_), .D(_8235__bF_buf4), .Y(_8237_) );
	NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_8237_), .Y(_6735__1_) );
	AOI22X1 AOI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr1_2_), .D(_8235__bF_buf3), .Y(_8238_) );
	NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_8238_), .Y(_6735__2_) );
	AOI22X1 AOI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8233__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr1_3_), .D(_8235__bF_buf2), .Y(_8239_) );
	NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_8239_), .Y(_6735__3_) );
	AOI22X1 AOI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr1_4_), .D(_8235__bF_buf1), .Y(_8240_) );
	NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf70), .B(_8240_), .Y(_6735__4_) );
	AOI22X1 AOI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8233__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr1_5_), .D(_8235__bF_buf0), .Y(_8241_) );
	NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf69), .B(_8241_), .Y(_6735__5_) );
	AOI22X1 AOI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8233__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr1_6_), .D(_8235__bF_buf5), .Y(_8242_) );
	NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_8242_), .Y(_6735__6_) );
	AOI22X1 AOI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr1_7_), .D(_8235__bF_buf4), .Y(_8243_) );
	NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf67), .B(_8243_), .Y(_6735__7_) );
	AOI22X1 AOI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr1_8_), .D(_8235__bF_buf3), .Y(_8244_) );
	NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf66), .B(_8244_), .Y(_6735__8_) );
	AOI22X1 AOI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8233__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr1_9_), .D(_8235__bF_buf2), .Y(_8245_) );
	NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf65), .B(_8245_), .Y(_6735__9_) );
	AOI22X1 AOI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr1_10_), .D(_8235__bF_buf1), .Y(_8246_) );
	NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf64), .B(_8246_), .Y(_6735__10_) );
	AOI22X1 AOI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8233__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr1_11_), .D(_8235__bF_buf0), .Y(_8247_) );
	NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf63), .B(_8247_), .Y(_6735__11_) );
	AOI22X1 AOI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8233__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr1_12_), .D(_8235__bF_buf5), .Y(_8248_) );
	NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf62), .B(_8248_), .Y(_6735__12_) );
	INVX1 INVX1_1412 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_13_), .Y(_8249_) );
	OAI21X1 OAI21X1_3514 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf2), .B(_8235__bF_buf4), .C(_6879__bF_buf6), .Y(_8250_) );
	AOI21X1 AOI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_8249_), .B(_8235__bF_buf3), .C(_8250_), .Y(_6735__13_) );
	AOI22X1 AOI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr1_14_), .D(_8235__bF_buf2), .Y(_8251_) );
	NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf61), .B(_8251_), .Y(_6735__14_) );
	INVX1 INVX1_1413 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_15_), .Y(_8252_) );
	OAI21X1 OAI21X1_3515 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf3), .B(_8235__bF_buf1), .C(_6879__bF_buf5), .Y(_8253_) );
	AOI21X1 AOI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_8252_), .B(_8235__bF_buf0), .C(_8253_), .Y(_6735__15_) );
	AOI22X1 AOI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr1_16_), .D(_8235__bF_buf5), .Y(_8254_) );
	NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf60), .B(_8254_), .Y(_6735__16_) );
	INVX1 INVX1_1414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_17_), .Y(_8255_) );
	OAI21X1 OAI21X1_3516 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf0), .B(_8235__bF_buf4), .C(_6879__bF_buf4), .Y(_8256_) );
	AOI21X1 AOI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_8255_), .B(_8235__bF_buf3), .C(_8256_), .Y(_6735__17_) );
	AOI22X1 AOI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8233__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr1_18_), .D(_8235__bF_buf2), .Y(_8257_) );
	NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf59), .B(_8257_), .Y(_6735__18_) );
	INVX1 INVX1_1415 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_19_), .Y(_8258_) );
	OAI21X1 OAI21X1_3517 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf1), .B(_8235__bF_buf1), .C(_6879__bF_buf3), .Y(_8259_) );
	AOI21X1 AOI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_8258_), .B(_8235__bF_buf0), .C(_8259_), .Y(_6735__19_) );
	AOI22X1 AOI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr1_20_), .D(_8235__bF_buf5), .Y(_8260_) );
	NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf58), .B(_8260_), .Y(_6735__20_) );
	INVX1 INVX1_1416 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_21_), .Y(_8261_) );
	OAI21X1 OAI21X1_3518 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf1), .B(_8235__bF_buf4), .C(_6879__bF_buf2), .Y(_8262_) );
	AOI21X1 AOI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_8261_), .B(_8235__bF_buf3), .C(_8262_), .Y(_6735__21_) );
	AOI22X1 AOI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8233__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr1_22_), .D(_8235__bF_buf2), .Y(_8263_) );
	NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf57), .B(_8263_), .Y(_6735__22_) );
	INVX1 INVX1_1417 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_23_), .Y(_8264_) );
	OAI21X1 OAI21X1_3519 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf3), .B(_8235__bF_buf1), .C(_6879__bF_buf1), .Y(_8265_) );
	AOI21X1 AOI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_8264_), .B(_8235__bF_buf0), .C(_8265_), .Y(_6735__23_) );
	AOI22X1 AOI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_8233__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr1_24_), .D(_8235__bF_buf5), .Y(_8266_) );
	NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf56), .B(_8266_), .Y(_6735__24_) );
	INVX1 INVX1_1418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_25_), .Y(_8267_) );
	OAI21X1 OAI21X1_3520 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf1), .B(_8235__bF_buf4), .C(_6879__bF_buf0), .Y(_8268_) );
	AOI21X1 AOI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(_8235__bF_buf3), .C(_8268_), .Y(_6735__25_) );
	AOI22X1 AOI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(_7406_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr1_26_), .D(_8235__bF_buf2), .Y(_8269_) );
	NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf55), .B(_8269_), .Y(_6735__26_) );
	INVX1 INVX1_1419 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_27_), .Y(_8270_) );
	OAI21X1 OAI21X1_3521 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf1), .B(_8235__bF_buf1), .C(_6879__bF_buf42), .Y(_8271_) );
	AOI21X1 AOI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_8270_), .B(_8235__bF_buf0), .C(_8271_), .Y(_6735__27_) );
	AOI22X1 AOI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr1_28_), .D(_8235__bF_buf5), .Y(_8272_) );
	NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf54), .B(_8272_), .Y(_6735__28_) );
	INVX1 INVX1_1420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_29_), .Y(_8273_) );
	OAI21X1 OAI21X1_3522 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf1), .B(_8235__bF_buf4), .C(_6879__bF_buf41), .Y(_8274_) );
	AOI21X1 AOI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .B(_8235__bF_buf3), .C(_8274_), .Y(_6735__29_) );
	AOI22X1 AOI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8233__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr1_30_), .D(_8235__bF_buf2), .Y(_8275_) );
	NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf53), .B(_8275_), .Y(_6735__30_) );
	INVX1 INVX1_1421 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_31_), .Y(_8276_) );
	OAI21X1 OAI21X1_3523 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf3), .B(_8235__bF_buf1), .C(_6879__bF_buf40), .Y(_8277_) );
	AOI21X1 AOI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_8276_), .B(_8235__bF_buf0), .C(_8277_), .Y(_6735__31_) );
	NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_8111__bF_buf2), .Y(_8278_) );
	NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_8278_), .Y(_8279_) );
	INVX8 INVX8_71 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .Y(_8280_) );
	NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8_bF_buf1), .B(_8280__bF_buf5), .Y(_8281_) );
	AOI22X1 AOI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8280__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr0_0_), .D(_8281__bF_buf5), .Y(_8282_) );
	NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf52), .B(_8282_), .Y(_6734__0_) );
	AOI22X1 AOI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8280__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_1_), .D(_8281__bF_buf4), .Y(_8283_) );
	NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf51), .B(_8283_), .Y(_6734__1_) );
	AOI22X1 AOI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8280__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_2_), .D(_8281__bF_buf3), .Y(_8284_) );
	NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf50), .B(_8284_), .Y(_6734__2_) );
	AOI22X1 AOI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8280__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr0_3_), .D(_8281__bF_buf2), .Y(_8285_) );
	NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf49), .B(_8285_), .Y(_6734__3_) );
	AOI22X1 AOI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8280__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr0_4_), .D(_8281__bF_buf1), .Y(_8286_) );
	NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf48), .B(_8286_), .Y(_6734__4_) );
	AOI22X1 AOI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8280__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr0_5_), .D(_8281__bF_buf0), .Y(_8287_) );
	NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf47), .B(_8287_), .Y(_6734__5_) );
	AOI22X1 AOI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8280__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr0_6_), .D(_8281__bF_buf5), .Y(_8288_) );
	NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf46), .B(_8288_), .Y(_6734__6_) );
	AOI22X1 AOI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8280__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_7_), .D(_8281__bF_buf4), .Y(_8289_) );
	NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf45), .B(_8289_), .Y(_6734__7_) );
	AOI22X1 AOI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8280__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_8_), .D(_8281__bF_buf3), .Y(_8290_) );
	NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf44), .B(_8290_), .Y(_6734__8_) );
	AOI22X1 AOI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8280__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr0_9_), .D(_8281__bF_buf2), .Y(_8291_) );
	NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf43), .B(_8291_), .Y(_6734__9_) );
	AOI22X1 AOI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8280__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr0_10_), .D(_8281__bF_buf1), .Y(_8292_) );
	NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf42), .B(_8292_), .Y(_6734__10_) );
	AOI22X1 AOI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8280__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr0_11_), .D(_8281__bF_buf0), .Y(_8293_) );
	NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf41), .B(_8293_), .Y(_6734__11_) );
	AOI22X1 AOI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8280__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr0_12_), .D(_8281__bF_buf5), .Y(_8294_) );
	NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf40), .B(_8294_), .Y(_6734__12_) );
	INVX1 INVX1_1422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_13_), .Y(_8295_) );
	OAI21X1 OAI21X1_3524 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf1), .B(_8281__bF_buf4), .C(_6879__bF_buf39), .Y(_8296_) );
	AOI21X1 AOI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_8295_), .B(_8281__bF_buf3), .C(_8296_), .Y(_6734__13_) );
	AOI22X1 AOI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8280__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_14_), .D(_8281__bF_buf2), .Y(_8297_) );
	NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf39), .B(_8297_), .Y(_6734__14_) );
	INVX1 INVX1_1423 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_15_), .Y(_8298_) );
	OAI21X1 OAI21X1_3525 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf2), .B(_8281__bF_buf1), .C(_6879__bF_buf38), .Y(_8299_) );
	AOI21X1 AOI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8281__bF_buf0), .C(_8299_), .Y(_6734__15_) );
	AOI22X1 AOI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_8280__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_16_), .D(_8281__bF_buf5), .Y(_8300_) );
	NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf38), .B(_8300_), .Y(_6734__16_) );
	INVX1 INVX1_1424 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_17_), .Y(_8301_) );
	OAI21X1 OAI21X1_3526 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf3), .B(_8281__bF_buf4), .C(_6879__bF_buf37), .Y(_8302_) );
	AOI21X1 AOI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_8301_), .B(_8281__bF_buf3), .C(_8302_), .Y(_6734__17_) );
	AOI22X1 AOI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8280__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr0_18_), .D(_8281__bF_buf2), .Y(_8303_) );
	NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf37), .B(_8303_), .Y(_6734__18_) );
	INVX1 INVX1_1425 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_19_), .Y(_8304_) );
	OAI21X1 OAI21X1_3527 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf0), .B(_8281__bF_buf1), .C(_6879__bF_buf36), .Y(_8305_) );
	AOI21X1 AOI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_8304_), .B(_8281__bF_buf0), .C(_8305_), .Y(_6734__19_) );
	AOI22X1 AOI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8280__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr0_20_), .D(_8281__bF_buf5), .Y(_8306_) );
	NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf36), .B(_8306_), .Y(_6734__20_) );
	INVX1 INVX1_1426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_21_), .Y(_8307_) );
	OAI21X1 OAI21X1_3528 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf0), .B(_8281__bF_buf4), .C(_6879__bF_buf35), .Y(_8308_) );
	AOI21X1 AOI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_8307_), .B(_8281__bF_buf3), .C(_8308_), .Y(_6734__21_) );
	AOI22X1 AOI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8280__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr0_22_), .D(_8281__bF_buf2), .Y(_8309_) );
	NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf35), .B(_8309_), .Y(_6734__22_) );
	INVX1 INVX1_1427 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_23_), .Y(_8310_) );
	OAI21X1 OAI21X1_3529 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf2), .B(_8281__bF_buf1), .C(_6879__bF_buf34), .Y(_8311_) );
	AOI21X1 AOI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8281__bF_buf0), .C(_8311_), .Y(_6734__23_) );
	AOI22X1 AOI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_8280__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr0_24_), .D(_8281__bF_buf5), .Y(_8312_) );
	NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf34), .B(_8312_), .Y(_6734__24_) );
	INVX1 INVX1_1428 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_25_), .Y(_8313_) );
	OAI21X1 OAI21X1_3530 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf0), .B(_8281__bF_buf4), .C(_6879__bF_buf33), .Y(_8314_) );
	AOI21X1 AOI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_8313_), .B(_8281__bF_buf3), .C(_8314_), .Y(_6734__25_) );
	AOI22X1 AOI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(_7406_), .B(_8280__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_26_), .D(_8281__bF_buf2), .Y(_8315_) );
	NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf33), .B(_8315_), .Y(_6734__26_) );
	INVX1 INVX1_1429 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_27_), .Y(_8316_) );
	OAI21X1 OAI21X1_3531 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf0), .B(_8281__bF_buf1), .C(_6879__bF_buf32), .Y(_8317_) );
	AOI21X1 AOI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_8316_), .B(_8281__bF_buf0), .C(_8317_), .Y(_6734__27_) );
	AOI22X1 AOI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8280__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_28_), .D(_8281__bF_buf5), .Y(_8318_) );
	NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf32), .B(_8318_), .Y(_6734__28_) );
	INVX1 INVX1_1430 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_29_), .Y(_8319_) );
	OAI21X1 OAI21X1_3532 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf0), .B(_8281__bF_buf4), .C(_6879__bF_buf31), .Y(_8320_) );
	AOI21X1 AOI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_8319_), .B(_8281__bF_buf3), .C(_8320_), .Y(_6734__29_) );
	AOI22X1 AOI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8280__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr0_30_), .D(_8281__bF_buf2), .Y(_8321_) );
	NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf31), .B(_8321_), .Y(_6734__30_) );
	INVX1 INVX1_1431 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_31_), .Y(_8322_) );
	OAI21X1 OAI21X1_3533 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf2), .B(_8281__bF_buf1), .C(_6879__bF_buf30), .Y(_8323_) );
	AOI21X1 AOI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(_8281__bF_buf0), .C(_8323_), .Y(_6734__31_) );
	NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf2), .B(_8113_), .Y(_8324_) );
	NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .B(_8324_), .Y(_8325_) );
	NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(_8231_), .Y(_8326_) );
	INVX8 INVX8_72 ( .gnd(gnd), .vdd(vdd), .A(_8326_), .Y(_8327_) );
	NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7_bF_buf1), .B(_8327__bF_buf6), .Y(_8328_) );
	AOI22X1 AOI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_8327__bF_buf5), .C(csr_gpr_iu_csr_pmp7cfg_0_), .D(_8328__bF_buf5), .Y(_8329_) );
	NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf30), .B(_8329_), .Y(_6733__0_) );
	INVX1 INVX1_1432 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_1_), .Y(_8330_) );
	OAI21X1 OAI21X1_3534 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_8328__bF_buf4), .C(_6879__bF_buf29), .Y(_8331_) );
	AOI21X1 AOI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_8330_), .B(_8328__bF_buf3), .C(_8331_), .Y(_6733__1_) );
	AOI22X1 AOI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(_7406_), .B(_8327__bF_buf4), .C(csr_gpr_iu_csr_pmp7cfg_2_), .D(_8328__bF_buf2), .Y(_8332_) );
	NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf29), .B(_8332_), .Y(_6733__2_) );
	INVX1 INVX1_1433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_3_), .Y(_8333_) );
	OAI21X1 OAI21X1_3535 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_8328__bF_buf1), .C(_6879__bF_buf28), .Y(_8334_) );
	AOI21X1 AOI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_8333_), .B(_8328__bF_buf0), .C(_8334_), .Y(_6733__3_) );
	AOI22X1 AOI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmp7cfg_4_), .D(_8328__bF_buf5), .Y(_8335_) );
	NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf28), .B(_8335_), .Y(_6733__4_) );
	INVX1 INVX1_1434 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_5_), .Y(_8336_) );
	OAI21X1 OAI21X1_3536 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_8328__bF_buf4), .C(_6879__bF_buf27), .Y(_8337_) );
	AOI21X1 AOI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_8336_), .B(_8328__bF_buf3), .C(_8337_), .Y(_6733__5_) );
	AOI22X1 AOI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmp7cfg_6_), .D(_8328__bF_buf2), .Y(_8338_) );
	NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf27), .B(_8338_), .Y(_6733__6_) );
	INVX1 INVX1_1435 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_7_), .Y(_8339_) );
	OAI21X1 OAI21X1_3537 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf1), .B(_8328__bF_buf1), .C(_6879__bF_buf26), .Y(_8340_) );
	AOI21X1 AOI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_8339_), .B(_8328__bF_buf0), .C(_8340_), .Y(_6733__7_) );
	AOI22X1 AOI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_8327__bF_buf1), .C(csr_gpr_iu_csr_pmp6cfg_0_), .D(_8328__bF_buf5), .Y(_8341_) );
	NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf26), .B(_8341_), .Y(_6732__0_) );
	INVX1 INVX1_1436 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_1_), .Y(_8342_) );
	OAI21X1 OAI21X1_3538 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf2), .B(_8328__bF_buf4), .C(_6879__bF_buf25), .Y(_8343_) );
	AOI21X1 AOI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_8342_), .B(_8328__bF_buf3), .C(_8343_), .Y(_6732__1_) );
	AOI22X1 AOI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_pmp6cfg_2_), .D(_8328__bF_buf2), .Y(_8344_) );
	NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf25), .B(_8344_), .Y(_6732__2_) );
	INVX1 INVX1_1437 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_3_), .Y(_8345_) );
	OAI21X1 OAI21X1_3539 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_8328__bF_buf1), .C(_6879__bF_buf24), .Y(_8346_) );
	AOI21X1 AOI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_8345_), .B(_8328__bF_buf0), .C(_8346_), .Y(_6732__3_) );
	AOI22X1 AOI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8327__bF_buf6), .C(csr_gpr_iu_csr_pmp6cfg_4_), .D(_8328__bF_buf5), .Y(_8347_) );
	NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf24), .B(_8347_), .Y(_6732__4_) );
	INVX1 INVX1_1438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_5_), .Y(_8348_) );
	OAI21X1 OAI21X1_3540 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_8328__bF_buf4), .C(_6879__bF_buf23), .Y(_8349_) );
	AOI21X1 AOI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_8348_), .B(_8328__bF_buf3), .C(_8349_), .Y(_6732__5_) );
	AOI22X1 AOI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8327__bF_buf5), .C(csr_gpr_iu_csr_pmp6cfg_6_), .D(_8328__bF_buf2), .Y(_8350_) );
	NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf23), .B(_8350_), .Y(_6732__6_) );
	INVX1 INVX1_1439 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_7_), .Y(_8351_) );
	OAI21X1 OAI21X1_3541 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf1), .B(_8328__bF_buf1), .C(_6879__bF_buf22), .Y(_8352_) );
	AOI21X1 AOI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_8351_), .B(_8328__bF_buf0), .C(_8352_), .Y(_6732__7_) );
	AOI22X1 AOI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8327__bF_buf4), .C(csr_gpr_iu_csr_pmp5cfg_0_), .D(_8328__bF_buf5), .Y(_8353_) );
	NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf22), .B(_8353_), .Y(_6731__0_) );
	AOI22X1 AOI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmp5cfg_1_), .D(_8328__bF_buf4), .Y(_8354_) );
	NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf21), .B(_8354_), .Y(_6731__1_) );
	AOI22X1 AOI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmp5cfg_2_), .D(_8328__bF_buf3), .Y(_8355_) );
	NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf20), .B(_8355_), .Y(_6731__2_) );
	AOI22X1 AOI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8327__bF_buf1), .C(csr_gpr_iu_csr_pmp5cfg_3_), .D(_8328__bF_buf2), .Y(_8356_) );
	NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf19), .B(_8356_), .Y(_6731__3_) );
	AOI22X1 AOI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_pmp5cfg_4_), .D(_8328__bF_buf1), .Y(_8357_) );
	NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf18), .B(_8357_), .Y(_6731__4_) );
	INVX1 INVX1_1440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_5_), .Y(_8358_) );
	OAI21X1 OAI21X1_3542 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf0), .B(_8328__bF_buf0), .C(_6879__bF_buf21), .Y(_8359_) );
	AOI21X1 AOI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_8358_), .B(_8328__bF_buf5), .C(_8359_), .Y(_6731__5_) );
	AOI22X1 AOI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8327__bF_buf6), .C(csr_gpr_iu_csr_pmp5cfg_6_), .D(_8328__bF_buf4), .Y(_8360_) );
	NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf17), .B(_8360_), .Y(_6731__6_) );
	INVX1 INVX1_1441 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_7_), .Y(_8361_) );
	OAI21X1 OAI21X1_3543 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf1), .B(_8328__bF_buf3), .C(_6879__bF_buf20), .Y(_8362_) );
	AOI21X1 AOI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_8361_), .B(_8328__bF_buf2), .C(_8362_), .Y(_6731__7_) );
	AOI22X1 AOI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8327__bF_buf5), .C(csr_gpr_iu_csr_pmp4cfg_0_), .D(_8328__bF_buf1), .Y(_8363_) );
	NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf16), .B(_8363_), .Y(_6730__0_) );
	AOI22X1 AOI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8327__bF_buf4), .C(csr_gpr_iu_csr_pmp4cfg_1_), .D(_8328__bF_buf0), .Y(_8364_) );
	NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf15), .B(_8364_), .Y(_6730__1_) );
	AOI22X1 AOI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmp4cfg_2_), .D(_8328__bF_buf5), .Y(_8365_) );
	NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf14), .B(_8365_), .Y(_6730__2_) );
	AOI22X1 AOI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmp4cfg_3_), .D(_8328__bF_buf4), .Y(_8366_) );
	NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf13), .B(_8366_), .Y(_6730__3_) );
	AOI22X1 AOI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8327__bF_buf1), .C(csr_gpr_iu_csr_pmp4cfg_4_), .D(_8328__bF_buf3), .Y(_8367_) );
	NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf12), .B(_8367_), .Y(_6730__4_) );
	AOI22X1 AOI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_pmp4cfg_5_), .D(_8328__bF_buf2), .Y(_8368_) );
	NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf11), .B(_8368_), .Y(_6730__5_) );
	AOI22X1 AOI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8327__bF_buf6), .C(csr_gpr_iu_csr_pmp4cfg_6_), .D(_8328__bF_buf1), .Y(_8369_) );
	NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf10), .B(_8369_), .Y(_6730__6_) );
	AOI22X1 AOI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8327__bF_buf5), .C(csr_gpr_iu_csr_pmp4cfg_7_), .D(_8328__bF_buf0), .Y(_8370_) );
	NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf9), .B(_8370_), .Y(_6730__7_) );
	NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(_8278_), .Y(_8371_) );
	INVX8 INVX8_73 ( .gnd(gnd), .vdd(vdd), .A(_8371_), .Y(_8372_) );
	NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6_bF_buf1), .B(_8372__bF_buf6), .Y(_8373_) );
	AOI22X1 AOI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_8372__bF_buf5), .C(csr_gpr_iu_csr_pmp3cfg_0_), .D(_8373__bF_buf5), .Y(_8374_) );
	NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf8), .B(_8374_), .Y(_6729__0_) );
	INVX1 INVX1_1442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp3cfg_1_), .Y(_8375_) );
	OAI21X1 OAI21X1_3544 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf2), .B(_8373__bF_buf4), .C(_6879__bF_buf19), .Y(_8376_) );
	AOI21X1 AOI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_8375_), .B(_8373__bF_buf3), .C(_8376_), .Y(_6729__1_) );
	AOI22X1 AOI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(_7406_), .B(_8372__bF_buf4), .C(csr_gpr_iu_csr_pmp3cfg_2_), .D(_8373__bF_buf2), .Y(_8377_) );
	NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf7), .B(_8377_), .Y(_6729__2_) );
	INVX1 INVX1_1443 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp3cfg_3_), .Y(_8378_) );
	OAI21X1 OAI21X1_3545 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf2), .B(_8373__bF_buf1), .C(_6879__bF_buf18), .Y(_8379_) );
	AOI21X1 AOI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_8378_), .B(_8373__bF_buf0), .C(_8379_), .Y(_6729__3_) );
	AOI22X1 AOI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8372__bF_buf3), .C(csr_gpr_iu_csr_pmp3cfg_4_), .D(_8373__bF_buf5), .Y(_8380_) );
	NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf6), .B(_8380_), .Y(_6729__4_) );
	INVX1 INVX1_1444 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp3cfg_5_), .Y(_8381_) );
	OAI21X1 OAI21X1_3546 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf2), .B(_8373__bF_buf4), .C(_6879__bF_buf17), .Y(_8382_) );
	AOI21X1 AOI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_8381_), .B(_8373__bF_buf3), .C(_8382_), .Y(_6729__5_) );
	AOI22X1 AOI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8372__bF_buf2), .C(csr_gpr_iu_csr_pmp3cfg_6_), .D(_8373__bF_buf2), .Y(_8383_) );
	NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .B(_8383_), .Y(_6729__6_) );
	INVX1 INVX1_1445 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp3cfg_7_), .Y(_8384_) );
	OAI21X1 OAI21X1_3547 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf0), .B(_8373__bF_buf1), .C(_6879__bF_buf16), .Y(_8385_) );
	AOI21X1 AOI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_8384_), .B(_8373__bF_buf0), .C(_8385_), .Y(_6729__7_) );
	AOI22X1 AOI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_8372__bF_buf1), .C(csr_gpr_iu_csr_pmp2cfg_0_), .D(_8373__bF_buf5), .Y(_8386_) );
	NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_8386_), .Y(_6728__0_) );
	INVX1 INVX1_1446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp2cfg_1_), .Y(_8387_) );
	OAI21X1 OAI21X1_3548 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf1), .B(_8373__bF_buf4), .C(_6879__bF_buf15), .Y(_8388_) );
	AOI21X1 AOI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_8387_), .B(_8373__bF_buf3), .C(_8388_), .Y(_6728__1_) );
	AOI22X1 AOI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8372__bF_buf0), .C(csr_gpr_iu_csr_pmp2cfg_2_), .D(_8373__bF_buf2), .Y(_8389_) );
	NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_8389_), .Y(_6728__2_) );
	INVX1 INVX1_1447 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp2cfg_3_), .Y(_8390_) );
	OAI21X1 OAI21X1_3549 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf2), .B(_8373__bF_buf1), .C(_6879__bF_buf14), .Y(_8391_) );
	AOI21X1 AOI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_8390_), .B(_8373__bF_buf0), .C(_8391_), .Y(_6728__3_) );
	AOI22X1 AOI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8372__bF_buf6), .C(csr_gpr_iu_csr_pmp2cfg_4_), .D(_8373__bF_buf5), .Y(_8392_) );
	NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_8392_), .Y(_6728__4_) );
	INVX1 INVX1_1448 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp2cfg_5_), .Y(_8393_) );
	OAI21X1 OAI21X1_3550 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf2), .B(_8373__bF_buf4), .C(_6879__bF_buf13), .Y(_8394_) );
	AOI21X1 AOI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_8393_), .B(_8373__bF_buf3), .C(_8394_), .Y(_6728__5_) );
	AOI22X1 AOI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8372__bF_buf5), .C(csr_gpr_iu_csr_pmp2cfg_6_), .D(_8373__bF_buf2), .Y(_8395_) );
	NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_8395_), .Y(_6728__6_) );
	INVX1 INVX1_1449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp2cfg_7_), .Y(_8396_) );
	OAI21X1 OAI21X1_3551 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf0), .B(_8373__bF_buf1), .C(_6879__bF_buf12), .Y(_8397_) );
	AOI21X1 AOI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_8396_), .B(_8373__bF_buf0), .C(_8397_), .Y(_6728__7_) );
	AOI22X1 AOI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8372__bF_buf4), .C(csr_gpr_iu_csr_pmp1cfg_0_), .D(_8373__bF_buf5), .Y(_8398_) );
	NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_8398_), .Y(_6727__0_) );
	AOI22X1 AOI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8372__bF_buf3), .C(csr_gpr_iu_csr_pmp1cfg_1_), .D(_8373__bF_buf4), .Y(_8399_) );
	NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf70), .B(_8399_), .Y(_6727__1_) );
	AOI22X1 AOI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8372__bF_buf2), .C(csr_gpr_iu_csr_pmp1cfg_2_), .D(_8373__bF_buf3), .Y(_8400_) );
	NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf69), .B(_8400_), .Y(_6727__2_) );
	AOI22X1 AOI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8372__bF_buf1), .C(csr_gpr_iu_csr_pmp1cfg_3_), .D(_8373__bF_buf2), .Y(_8401_) );
	NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_8401_), .Y(_6727__3_) );
	AOI22X1 AOI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8372__bF_buf0), .C(csr_gpr_iu_csr_pmp1cfg_4_), .D(_8373__bF_buf1), .Y(_8402_) );
	NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf67), .B(_8402_), .Y(_6727__4_) );
	INVX1 INVX1_1450 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp1cfg_5_), .Y(_8403_) );
	OAI21X1 OAI21X1_3552 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_8373__bF_buf0), .C(_6879__bF_buf11), .Y(_8404_) );
	AOI21X1 AOI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_8403_), .B(_8373__bF_buf5), .C(_8404_), .Y(_6727__5_) );
	AOI22X1 AOI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8372__bF_buf6), .C(csr_gpr_iu_csr_pmp1cfg_6_), .D(_8373__bF_buf4), .Y(_8405_) );
	NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf66), .B(_8405_), .Y(_6727__6_) );
	INVX1 INVX1_1451 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp1cfg_7_), .Y(_8406_) );
	OAI21X1 OAI21X1_3553 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf0), .B(_8373__bF_buf3), .C(_6879__bF_buf10), .Y(_8407_) );
	AOI21X1 AOI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_8406_), .B(_8373__bF_buf2), .C(_8407_), .Y(_6727__7_) );
	AOI22X1 AOI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8372__bF_buf5), .C(csr_gpr_iu_csr_pmp0cfg_0_), .D(_8373__bF_buf1), .Y(_8408_) );
	NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf65), .B(_8408_), .Y(_6726__0_) );
	AOI22X1 AOI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8372__bF_buf4), .C(csr_gpr_iu_csr_pmp0cfg_1_), .D(_8373__bF_buf0), .Y(_8409_) );
	NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf64), .B(_8409_), .Y(_6726__1_) );
	AOI22X1 AOI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8372__bF_buf3), .C(csr_gpr_iu_csr_pmp0cfg_2_), .D(_8373__bF_buf5), .Y(_8410_) );
	NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf63), .B(_8410_), .Y(_6726__2_) );
	AOI22X1 AOI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8372__bF_buf2), .C(csr_gpr_iu_csr_pmp0cfg_3_), .D(_8373__bF_buf4), .Y(_8411_) );
	NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf62), .B(_8411_), .Y(_6726__3_) );
	AOI22X1 AOI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8372__bF_buf1), .C(csr_gpr_iu_csr_pmp0cfg_4_), .D(_8373__bF_buf3), .Y(_8412_) );
	NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf61), .B(_8412_), .Y(_6726__4_) );
	AOI22X1 AOI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8372__bF_buf0), .C(csr_gpr_iu_csr_pmp0cfg_5_), .D(_8373__bF_buf2), .Y(_8413_) );
	NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf60), .B(_8413_), .Y(_6726__5_) );
	AOI22X1 AOI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8372__bF_buf6), .C(csr_gpr_iu_csr_pmp0cfg_6_), .D(_8373__bF_buf1), .Y(_8414_) );
	NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf59), .B(_8414_), .Y(_6726__6_) );
	AOI22X1 AOI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8372__bF_buf5), .C(csr_gpr_iu_csr_pmp0cfg_7_), .D(_8373__bF_buf0), .Y(_8415_) );
	NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf58), .B(_8415_), .Y(_6726__7_) );
	NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_8278_), .Y(_8416_) );
	INVX8 INVX8_74 ( .gnd(gnd), .vdd(vdd), .A(_8416_), .Y(_8417_) );
	NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_8416_), .Y(_8418_) );
	INVX8 INVX8_75 ( .gnd(gnd), .vdd(vdd), .A(_8418_), .Y(_8419_) );
	AOI22X1 AOI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8417__bF_buf5), .C(csr_gpr_iu_csr_mscratch_0_), .D(_8419__bF_buf5), .Y(_8420_) );
	NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf57), .B(_8420_), .Y(_6716__0_) );
	AOI22X1 AOI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8417__bF_buf4), .C(csr_gpr_iu_csr_mscratch_1_), .D(_8419__bF_buf4), .Y(_8421_) );
	NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf56), .B(_8421_), .Y(_6716__1_) );
	AOI22X1 AOI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8417__bF_buf3), .C(csr_gpr_iu_csr_mscratch_2_), .D(_8419__bF_buf3), .Y(_8422_) );
	NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf55), .B(_8422_), .Y(_6716__2_) );
	AOI22X1 AOI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8417__bF_buf2), .C(csr_gpr_iu_csr_mscratch_3_), .D(_8419__bF_buf2), .Y(_8423_) );
	NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf54), .B(_8423_), .Y(_6716__3_) );
	AOI22X1 AOI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8417__bF_buf1), .C(csr_gpr_iu_csr_mscratch_4_), .D(_8419__bF_buf1), .Y(_8424_) );
	NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf53), .B(_8424_), .Y(_6716__4_) );
	AOI22X1 AOI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8417__bF_buf0), .C(csr_gpr_iu_csr_mscratch_5_), .D(_8419__bF_buf0), .Y(_8425_) );
	NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf52), .B(_8425_), .Y(_6716__5_) );
	AOI22X1 AOI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8417__bF_buf5), .C(csr_gpr_iu_csr_mscratch_6_), .D(_8419__bF_buf5), .Y(_8426_) );
	NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf51), .B(_8426_), .Y(_6716__6_) );
	AOI22X1 AOI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8417__bF_buf4), .C(csr_gpr_iu_csr_mscratch_7_), .D(_8419__bF_buf4), .Y(_8427_) );
	NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf50), .B(_8427_), .Y(_6716__7_) );
	AOI22X1 AOI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8417__bF_buf3), .C(csr_gpr_iu_csr_mscratch_8_), .D(_8419__bF_buf3), .Y(_8428_) );
	NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf49), .B(_8428_), .Y(_6716__8_) );
	AOI22X1 AOI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8417__bF_buf2), .C(csr_gpr_iu_csr_mscratch_9_), .D(_8419__bF_buf2), .Y(_8429_) );
	NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf48), .B(_8429_), .Y(_6716__9_) );
	AOI22X1 AOI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_8417__bF_buf1), .C(csr_gpr_iu_csr_mscratch_10_), .D(_8419__bF_buf1), .Y(_8430_) );
	NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf47), .B(_8430_), .Y(_6716__10_) );
	AOI22X1 AOI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8417__bF_buf0), .C(csr_gpr_iu_csr_mscratch_11_), .D(_8419__bF_buf0), .Y(_8431_) );
	NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf46), .B(_8431_), .Y(_6716__11_) );
	AOI22X1 AOI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .B(_8417__bF_buf5), .C(csr_gpr_iu_csr_mscratch_12_), .D(_8419__bF_buf5), .Y(_8432_) );
	NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf45), .B(_8432_), .Y(_6716__12_) );
	INVX1 INVX1_1452 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_13_), .Y(_8433_) );
	OAI21X1 OAI21X1_3554 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf2), .B(_8419__bF_buf4), .C(_6879__bF_buf9), .Y(_8434_) );
	AOI21X1 AOI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_8433_), .B(_8419__bF_buf3), .C(_8434_), .Y(_6716__13_) );
	AOI22X1 AOI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_8417__bF_buf4), .C(csr_gpr_iu_csr_mscratch_14_), .D(_8419__bF_buf2), .Y(_8435_) );
	NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf44), .B(_8435_), .Y(_6716__14_) );
	INVX1 INVX1_1453 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_15_), .Y(_8436_) );
	OAI21X1 OAI21X1_3555 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf3), .B(_8419__bF_buf1), .C(_6879__bF_buf8), .Y(_8437_) );
	AOI21X1 AOI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_8436_), .B(_8419__bF_buf0), .C(_8437_), .Y(_6716__15_) );
	OAI21X1 OAI21X1_3556 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_8416_), .C(csr_gpr_iu_csr_mscratch_16_), .Y(_8438_) );
	OAI21X1 OAI21X1_3557 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_8419__bF_buf5), .C(_8438_), .Y(_8439_) );
	AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_8439_), .B(_6879__bF_buf7), .Y(_6716__16_) );
	INVX1 INVX1_1454 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_17_), .Y(_8440_) );
	OAI21X1 OAI21X1_3558 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf0), .B(_8419__bF_buf4), .C(_6879__bF_buf6), .Y(_8441_) );
	AOI21X1 AOI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_8440_), .B(_8419__bF_buf3), .C(_8441_), .Y(_6716__17_) );
	AOI22X1 AOI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_8417__bF_buf3), .C(csr_gpr_iu_csr_mscratch_18_), .D(_8419__bF_buf2), .Y(_8442_) );
	NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf43), .B(_8442_), .Y(_6716__18_) );
	INVX1 INVX1_1455 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_19_), .Y(_8443_) );
	OAI21X1 OAI21X1_3559 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf1), .B(_8419__bF_buf1), .C(_6879__bF_buf5), .Y(_8444_) );
	AOI21X1 AOI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_8443_), .B(_8419__bF_buf0), .C(_8444_), .Y(_6716__19_) );
	AOI22X1 AOI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_8417__bF_buf2), .C(csr_gpr_iu_csr_mscratch_20_), .D(_8419__bF_buf5), .Y(_8445_) );
	NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf42), .B(_8445_), .Y(_6716__20_) );
	INVX1 INVX1_1456 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_21_), .Y(_8446_) );
	OAI21X1 OAI21X1_3560 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf1), .B(_8419__bF_buf4), .C(_6879__bF_buf4), .Y(_8447_) );
	AOI21X1 AOI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_8446_), .B(_8419__bF_buf3), .C(_8447_), .Y(_6716__21_) );
	AOI22X1 AOI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_8417__bF_buf1), .C(csr_gpr_iu_csr_mscratch_22_), .D(_8419__bF_buf2), .Y(_8448_) );
	NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf41), .B(_8448_), .Y(_6716__22_) );
	INVX1 INVX1_1457 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_23_), .Y(_8449_) );
	OAI21X1 OAI21X1_3561 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf3), .B(_8419__bF_buf1), .C(_6879__bF_buf3), .Y(_8450_) );
	AOI21X1 AOI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_8449_), .B(_8419__bF_buf0), .C(_8450_), .Y(_6716__23_) );
	OAI21X1 OAI21X1_3562 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_8416_), .C(csr_gpr_iu_csr_mscratch_24_), .Y(_8451_) );
	OAI21X1 OAI21X1_3563 ( .gnd(gnd), .vdd(vdd), .A(_7399_), .B(_8419__bF_buf5), .C(_8451_), .Y(_8452_) );
	AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_8452_), .B(_6879__bF_buf2), .Y(_6716__24_) );
	INVX1 INVX1_1458 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_25_), .Y(_8453_) );
	OAI21X1 OAI21X1_3564 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf1), .B(_8419__bF_buf4), .C(_6879__bF_buf1), .Y(_8454_) );
	AOI21X1 AOI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_8453_), .B(_8419__bF_buf3), .C(_8454_), .Y(_6716__25_) );
	OAI21X1 OAI21X1_3565 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_8416_), .C(csr_gpr_iu_csr_mscratch_26_), .Y(_8455_) );
	OAI21X1 OAI21X1_3566 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_8419__bF_buf2), .C(_8455_), .Y(_8456_) );
	AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_8456_), .B(_6879__bF_buf0), .Y(_6716__26_) );
	INVX1 INVX1_1459 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_27_), .Y(_8457_) );
	OAI21X1 OAI21X1_3567 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf1), .B(_8419__bF_buf1), .C(_6879__bF_buf42), .Y(_8458_) );
	AOI21X1 AOI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_8457_), .B(_8419__bF_buf0), .C(_8458_), .Y(_6716__27_) );
	OAI21X1 OAI21X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_8416_), .C(csr_gpr_iu_csr_mscratch_28_), .Y(_8459_) );
	OAI21X1 OAI21X1_3569 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_8419__bF_buf5), .C(_8459_), .Y(_8460_) );
	AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_8460_), .B(_6879__bF_buf41), .Y(_6716__28_) );
	INVX1 INVX1_1460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_29_), .Y(_8461_) );
	OAI21X1 OAI21X1_3570 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf1), .B(_8419__bF_buf4), .C(_6879__bF_buf40), .Y(_8462_) );
	AOI21X1 AOI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_8461_), .B(_8419__bF_buf3), .C(_8462_), .Y(_6716__29_) );
	AOI22X1 AOI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(_7417_), .B(_8417__bF_buf0), .C(csr_gpr_iu_csr_mscratch_30_), .D(_8419__bF_buf2), .Y(_8463_) );
	NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf40), .B(_8463_), .Y(_6716__30_) );
	INVX1 INVX1_1461 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_31_), .Y(_8464_) );
	OAI21X1 OAI21X1_3571 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf3), .B(_8419__bF_buf1), .C(_6879__bF_buf39), .Y(_8465_) );
	AOI21X1 AOI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_8464_), .B(_8419__bF_buf0), .C(_8465_), .Y(_6716__31_) );
	NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_7311_), .B(_8058_), .Y(_8466_) );
	NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_8057_), .B(_8466_), .Y(_8467_) );
	INVX1 INVX1_1462 ( .gnd(gnd), .vdd(vdd), .A(_8467_), .Y(_8468_) );
	NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_8468_), .Y(_8469_) );
	INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .Y(_8470_) );
	OAI21X1 OAI21X1_3572 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(_8470_), .C(csr_gpr_iu_csr_ssie), .Y(_8471_) );
	NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_7329_), .Y(_8472_) );
	AOI21X1 AOI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_8471_), .B(_8472_), .C(rst_bF_buf39), .Y(_6747_) );
	NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_8107_), .B(_8470_), .Y(_8473_) );
	INVX1 INVX1_1463 ( .gnd(gnd), .vdd(vdd), .A(_8473_), .Y(_8474_) );
	OAI21X1 OAI21X1_3573 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf3), .B(_8474_), .C(csr_gpr_iu_csr_msie), .Y(_8475_) );
	NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8473_), .Y(_8476_) );
	AOI21X1 AOI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_8475_), .B(_8476_), .C(rst_bF_buf38), .Y(_6717_) );
	OAI21X1 OAI21X1_3574 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf3), .B(_8470_), .C(csr_gpr_iu_csr_stie), .Y(_8477_) );
	NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_7342_), .Y(_8478_) );
	AOI21X1 AOI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_8477_), .B(_8478_), .C(rst_bF_buf37), .Y(_6749_) );
	OAI21X1 OAI21X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf3), .B(_8474_), .C(csr_gpr_iu_csr_mtie), .Y(_8479_) );
	NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8473_), .Y(_8480_) );
	AOI21X1 AOI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_8479_), .B(_8480_), .C(rst_bF_buf36), .Y(_6720_) );
	OAI21X1 OAI21X1_3576 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf3), .B(_8470_), .C(csr_gpr_iu_csr_seie), .Y(_8481_) );
	NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_7303__bF_buf5_bF_buf1), .C(_8469_), .Y(_8482_) );
	AOI21X1 AOI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_8481_), .B(_8482_), .C(rst_bF_buf35), .Y(_6740_) );
	OAI21X1 OAI21X1_3577 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf3), .B(_8474_), .C(csr_gpr_iu_csr_meie), .Y(_8483_) );
	NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_8473_), .Y(_8484_) );
	AOI21X1 AOI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_8483_), .B(_8484_), .C(rst_bF_buf34), .Y(_6707_) );
	INVX1 INVX1_1464 ( .gnd(gnd), .vdd(vdd), .A(_8057_), .Y(_8485_) );
	NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_8485_), .B(_8161_), .Y(_8486_) );
	OAI21X1 OAI21X1_3578 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf3), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_0_), .Y(_8487_) );
	NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_8485_), .B(_7433_), .Y(_8488_) );
	NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_8488_), .Y(_8489_) );
	NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf5), .B(_7325_), .Y(_8490_) );
	AOI21X1 AOI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_8490_), .B(_8487_), .C(rst_bF_buf33), .Y(_6706__0_) );
	OAI21X1 OAI21X1_3579 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf3), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_1_), .Y(_8491_) );
	NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf4), .B(_7329_), .Y(_8492_) );
	AOI21X1 AOI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .B(_8491_), .C(rst_bF_buf32), .Y(_6706__1_) );
	OAI21X1 OAI21X1_3580 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf3), .B(_8486__bF_buf1), .C(csr_gpr_iu_csr_medeleg_2_), .Y(_8493_) );
	NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf3), .B(_7333_), .Y(_8494_) );
	AOI21X1 AOI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_8494_), .B(_8493_), .C(rst_bF_buf31), .Y(_6706__2_) );
	OAI21X1 OAI21X1_3581 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf3), .B(_8486__bF_buf0), .C(csr_gpr_iu_csr_medeleg_3_), .Y(_8495_) );
	NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf2), .B(_7336_), .Y(_8496_) );
	AOI21X1 AOI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_8496_), .B(_8495_), .C(rst_bF_buf30), .Y(_6706__3_) );
	OAI21X1 OAI21X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_4_), .Y(_8497_) );
	NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf1), .B(_7339_), .Y(_8498_) );
	AOI21X1 AOI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8497_), .C(rst_bF_buf29), .Y(_6706__4_) );
	OAI21X1 OAI21X1_3583 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_5_), .Y(_8499_) );
	NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf0), .B(_7342_), .Y(_8500_) );
	AOI21X1 AOI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_8500_), .B(_8499_), .C(rst_bF_buf28), .Y(_6706__5_) );
	OAI21X1 OAI21X1_3584 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_8486__bF_buf1), .C(csr_gpr_iu_csr_medeleg_6_), .Y(_8501_) );
	NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf5), .B(_7345_), .Y(_8502_) );
	AOI21X1 AOI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_8502_), .B(_8501_), .C(rst_bF_buf27), .Y(_6706__6_) );
	OAI21X1 OAI21X1_3585 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_8486__bF_buf0), .C(csr_gpr_iu_csr_medeleg_7_), .Y(_8503_) );
	NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf4), .B(_7348_), .Y(_8504_) );
	AOI21X1 AOI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_8504_), .B(_8503_), .C(rst_bF_buf26), .Y(_6706__7_) );
	OAI21X1 OAI21X1_3586 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_8_), .Y(_8505_) );
	NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf3), .B(_7351_), .Y(_8506_) );
	AOI21X1 AOI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_8506_), .B(_8505_), .C(rst_bF_buf25), .Y(_6706__8_) );
	OAI21X1 OAI21X1_3587 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_9_), .Y(_8507_) );
	NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf2), .B(_7354_), .Y(_8508_) );
	AOI21X1 AOI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_8508_), .B(_8507_), .C(rst_bF_buf24), .Y(_6706__9_) );
	OAI21X1 OAI21X1_3588 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf2), .B(_8486__bF_buf1), .C(csr_gpr_iu_csr_medeleg_10_), .Y(_8509_) );
	NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf1), .B(_7357_), .Y(_8510_) );
	AOI21X1 AOI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_8510_), .B(_8509_), .C(rst_bF_buf23), .Y(_6706__10_) );
	OAI21X1 OAI21X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf2), .B(_8486__bF_buf0), .C(csr_gpr_iu_csr_medeleg_11_), .Y(_8511_) );
	NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf0), .B(_7360_), .Y(_8512_) );
	AOI21X1 AOI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_8512_), .B(_8511_), .C(rst_bF_buf22), .Y(_6706__11_) );
	OAI21X1 OAI21X1_3590 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf2), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_12_), .Y(_8513_) );
	NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf5), .B(_7363_), .Y(_8514_) );
	AOI21X1 AOI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_8514_), .B(_8513_), .C(rst_bF_buf21), .Y(_6706__12_) );
	INVX1 INVX1_1465 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_13_), .Y(_8515_) );
	NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4_bF_buf1), .B(_8489__bF_buf4), .Y(_8516_) );
	OAI21X1 OAI21X1_3591 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf1), .B(_8516__bF_buf3), .C(_6879__bF_buf38), .Y(_8517_) );
	AOI21X1 AOI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_8515_), .B(_8516__bF_buf2), .C(_8517_), .Y(_6706__13_) );
	OAI21X1 OAI21X1_3592 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf2), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_14_), .Y(_8518_) );
	NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf3), .B(_7370_), .Y(_8519_) );
	AOI21X1 AOI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_8518_), .B(_8519_), .C(rst_bF_buf20), .Y(_6706__14_) );
	INVX1 INVX1_1466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_15_), .Y(_8520_) );
	OAI21X1 OAI21X1_3593 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf2), .B(_8516__bF_buf1), .C(_6879__bF_buf37), .Y(_8521_) );
	AOI21X1 AOI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_8520_), .B(_8516__bF_buf0), .C(_8521_), .Y(_6706__15_) );
	OAI21X1 OAI21X1_3594 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf2), .B(_8486__bF_buf1), .C(csr_gpr_iu_csr_medeleg_16_), .Y(_8522_) );
	NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf2), .B(_7376_), .Y(_8523_) );
	AOI21X1 AOI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_8522_), .B(_8523_), .C(rst_bF_buf19), .Y(_6706__16_) );
	INVX1 INVX1_1467 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_17_), .Y(_8524_) );
	OAI21X1 OAI21X1_3595 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf3), .B(_8516__bF_buf3), .C(_6879__bF_buf36), .Y(_8525_) );
	AOI21X1 AOI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_8524_), .B(_8516__bF_buf2), .C(_8525_), .Y(_6706__17_) );
	OAI21X1 OAI21X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf9_bF_buf2), .B(_8486__bF_buf0), .C(csr_gpr_iu_csr_medeleg_18_), .Y(_8526_) );
	NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf1), .B(_7382_), .Y(_8527_) );
	AOI21X1 AOI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_8526_), .B(_8527_), .C(rst_bF_buf18), .Y(_6706__18_) );
	INVX1 INVX1_1468 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_19_), .Y(_8528_) );
	OAI21X1 OAI21X1_3597 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf0), .B(_8516__bF_buf1), .C(_6879__bF_buf35), .Y(_8529_) );
	AOI21X1 AOI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_8528_), .B(_8516__bF_buf0), .C(_8529_), .Y(_6706__19_) );
	OAI21X1 OAI21X1_3598 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf8_bF_buf2), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_20_), .Y(_8530_) );
	NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf0), .B(_7388_), .Y(_8531_) );
	AOI21X1 AOI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_8530_), .B(_8531_), .C(rst_bF_buf17), .Y(_6706__20_) );
	INVX1 INVX1_1469 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_21_), .Y(_8532_) );
	OAI21X1 OAI21X1_3599 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf0), .B(_8516__bF_buf3), .C(_6879__bF_buf34), .Y(_8533_) );
	AOI21X1 AOI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_8532_), .B(_8516__bF_buf2), .C(_8533_), .Y(_6706__21_) );
	OAI21X1 OAI21X1_3600 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf7_bF_buf2), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_22_), .Y(_8534_) );
	NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf5), .B(_7394_), .Y(_8535_) );
	AOI21X1 AOI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_8534_), .B(_8535_), .C(rst_bF_buf16), .Y(_6706__22_) );
	INVX1 INVX1_1470 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_23_), .Y(_8536_) );
	OAI21X1 OAI21X1_3601 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf2), .B(_8516__bF_buf1), .C(_6879__bF_buf33), .Y(_8537_) );
	AOI21X1 AOI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_8536_), .B(_8516__bF_buf0), .C(_8537_), .Y(_6706__23_) );
	OAI21X1 OAI21X1_3602 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf6_bF_buf2), .B(_8486__bF_buf1), .C(csr_gpr_iu_csr_medeleg_24_), .Y(_8538_) );
	NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf4), .B(_7400_), .Y(_8539_) );
	AOI21X1 AOI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_8539_), .C(rst_bF_buf15), .Y(_6706__24_) );
	INVX1 INVX1_1471 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_25_), .Y(_8540_) );
	OAI21X1 OAI21X1_3603 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf0), .B(_8516__bF_buf3), .C(_6879__bF_buf32), .Y(_8541_) );
	AOI21X1 AOI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_8540_), .B(_8516__bF_buf2), .C(_8541_), .Y(_6706__25_) );
	OAI21X1 OAI21X1_3604 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf5), .B(_8486__bF_buf0), .C(csr_gpr_iu_csr_medeleg_26_), .Y(_8542_) );
	NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf3), .B(_7406_), .Y(_8543_) );
	AOI21X1 AOI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_8542_), .B(_8543_), .C(rst_bF_buf14), .Y(_6706__26_) );
	INVX1 INVX1_1472 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_27_), .Y(_8544_) );
	OAI21X1 OAI21X1_3605 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf0), .B(_8516__bF_buf1), .C(_6879__bF_buf31), .Y(_8545_) );
	AOI21X1 AOI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_8544_), .B(_8516__bF_buf0), .C(_8545_), .Y(_6706__27_) );
	OAI21X1 OAI21X1_3606 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf4), .B(_8486__bF_buf3), .C(csr_gpr_iu_csr_medeleg_28_), .Y(_8546_) );
	NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf2), .B(_7412_), .Y(_8547_) );
	AOI21X1 AOI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_8546_), .B(_8547_), .C(rst_bF_buf13), .Y(_6706__28_) );
	INVX1 INVX1_1473 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_29_), .Y(_8548_) );
	OAI21X1 OAI21X1_3607 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf0), .B(_8516__bF_buf3), .C(_6879__bF_buf30), .Y(_8549_) );
	AOI21X1 AOI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_8548_), .B(_8516__bF_buf2), .C(_8549_), .Y(_6706__29_) );
	OAI21X1 OAI21X1_3608 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf3), .B(_8486__bF_buf2), .C(csr_gpr_iu_csr_medeleg_30_), .Y(_8550_) );
	NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_8489__bF_buf1), .B(_7417_), .Y(_8551_) );
	AOI21X1 AOI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_8550_), .B(_8551_), .C(rst_bF_buf12), .Y(_6706__30_) );
	INVX1 INVX1_1474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_31_), .Y(_8552_) );
	OAI21X1 OAI21X1_3609 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf2), .B(_8516__bF_buf1), .C(_6879__bF_buf29), .Y(_8553_) );
	AOI21X1 AOI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_8552_), .B(_8516__bF_buf0), .C(_8553_), .Y(_6706__31_) );
	NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_8485_), .B(_8112_), .Y(_8554_) );
	INVX4 INVX4_18 ( .gnd(gnd), .vdd(vdd), .A(_8554_), .Y(_8555_) );
	NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_8554_), .Y(_8556_) );
	INVX8 INVX8_76 ( .gnd(gnd), .vdd(vdd), .A(_8556_), .Y(_8557_) );
	AOI22X1 AOI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_0_), .D(_8557__bF_buf5), .Y(_8558_) );
	NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf11), .B(_8558_), .Y(_6710__0_) );
	AOI22X1 AOI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_1_), .D(_8557__bF_buf4), .Y(_8559_) );
	NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf10), .B(_8559_), .Y(_6710__1_) );
	AOI22X1 AOI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_2_), .D(_8557__bF_buf3), .Y(_8560_) );
	NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf9), .B(_8560_), .Y(_6710__2_) );
	AOI22X1 AOI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_3_), .D(_8557__bF_buf2), .Y(_8561_) );
	NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf8), .B(_8561_), .Y(_6710__3_) );
	AOI22X1 AOI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_4_), .D(_8557__bF_buf1), .Y(_8562_) );
	NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf7), .B(_8562_), .Y(_6710__4_) );
	AOI22X1 AOI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_5_), .D(_8557__bF_buf0), .Y(_8563_) );
	NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf6), .B(_8563_), .Y(_6710__5_) );
	AOI22X1 AOI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_6_), .D(_8557__bF_buf5), .Y(_8564_) );
	NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .B(_8564_), .Y(_6710__6_) );
	AOI22X1 AOI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_7_), .D(_8557__bF_buf4), .Y(_8565_) );
	NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_8565_), .Y(_6710__7_) );
	AOI22X1 AOI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_8_), .D(_8557__bF_buf3), .Y(_8566_) );
	NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_8566_), .Y(_6710__8_) );
	AOI22X1 AOI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_8555_), .C(csr_gpr_iu_csr_mideleg_9_), .D(_8557__bF_buf2), .Y(_8567_) );
	NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_8567_), .Y(_6710__9_) );
	NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_8556_), .Y(_8568_) );
	OAI21X1 OAI21X1_3610 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_10_), .B(_8556_), .C(_8568_), .Y(_8569_) );
	NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_8569_), .Y(_6710__10_) );
	NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_8556_), .Y(_8570_) );
	OAI21X1 OAI21X1_3611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_11_), .B(_8556_), .C(_8570_), .Y(_8571_) );
	NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_8571_), .Y(_6710__11_) );
	OAI21X1 OAI21X1_3612 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_12_), .Y(_8572_) );
	OAI21X1 OAI21X1_3613 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_8557__bF_buf1), .C(_8572_), .Y(_8573_) );
	AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_8573_), .B(_6879__bF_buf28), .Y(_6710__12_) );
	INVX1 INVX1_1475 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_13_), .Y(_8574_) );
	OAI21X1 OAI21X1_3614 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf0), .B(_8557__bF_buf0), .C(_6879__bF_buf27), .Y(_8575_) );
	AOI21X1 AOI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_8574_), .B(_8557__bF_buf5), .C(_8575_), .Y(_6710__13_) );
	NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_8556_), .Y(_8576_) );
	OAI21X1 OAI21X1_3615 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_14_), .B(_8556_), .C(_8576_), .Y(_8577_) );
	NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf70), .B(_8577_), .Y(_6710__14_) );
	INVX1 INVX1_1476 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_15_), .Y(_8578_) );
	OAI21X1 OAI21X1_3616 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf1), .B(_8557__bF_buf4), .C(_6879__bF_buf26), .Y(_8579_) );
	AOI21X1 AOI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_8578_), .B(_8557__bF_buf3), .C(_8579_), .Y(_6710__15_) );
	OAI21X1 OAI21X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf0), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_16_), .Y(_8580_) );
	OAI21X1 OAI21X1_3618 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_8557__bF_buf2), .C(_8580_), .Y(_8581_) );
	AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_8581_), .B(_6879__bF_buf25), .Y(_6710__16_) );
	INVX1 INVX1_1477 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_17_), .Y(_8582_) );
	OAI21X1 OAI21X1_3619 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf2), .B(_8557__bF_buf1), .C(_6879__bF_buf24), .Y(_8583_) );
	AOI21X1 AOI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_8582_), .B(_8557__bF_buf0), .C(_8583_), .Y(_6710__17_) );
	NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_8556_), .Y(_8584_) );
	OAI21X1 OAI21X1_3620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_18_), .B(_8556_), .C(_8584_), .Y(_8585_) );
	NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf69), .B(_8585_), .Y(_6710__18_) );
	INVX1 INVX1_1478 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_19_), .Y(_8586_) );
	OAI21X1 OAI21X1_3621 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_8557__bF_buf5), .C(_6879__bF_buf23), .Y(_8587_) );
	AOI21X1 AOI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_8586_), .B(_8557__bF_buf4), .C(_8587_), .Y(_6710__19_) );
	OAI21X1 OAI21X1_3622 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf14_bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_20_), .Y(_8588_) );
	OAI21X1 OAI21X1_3623 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_8557__bF_buf3), .C(_8588_), .Y(_8589_) );
	AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_8589_), .B(_6879__bF_buf22), .Y(_6710__20_) );
	INVX1 INVX1_1479 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_21_), .Y(_8590_) );
	OAI21X1 OAI21X1_3624 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_8557__bF_buf2), .C(_6879__bF_buf21), .Y(_8591_) );
	AOI21X1 AOI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_8590_), .B(_8557__bF_buf1), .C(_8591_), .Y(_6710__21_) );
	OAI21X1 OAI21X1_3625 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf13_bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_22_), .Y(_8592_) );
	OAI21X1 OAI21X1_3626 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_8557__bF_buf0), .C(_8592_), .Y(_8593_) );
	AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_8593_), .B(_6879__bF_buf20), .Y(_6710__22_) );
	INVX1 INVX1_1480 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_23_), .Y(_8594_) );
	OAI21X1 OAI21X1_3627 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf1), .B(_8557__bF_buf5), .C(_6879__bF_buf19), .Y(_8595_) );
	AOI21X1 AOI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_8594_), .B(_8557__bF_buf4), .C(_8595_), .Y(_6710__23_) );
	OAI21X1 OAI21X1_3628 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf12_bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_24_), .Y(_8596_) );
	OAI21X1 OAI21X1_3629 ( .gnd(gnd), .vdd(vdd), .A(_7399_), .B(_8557__bF_buf3), .C(_8596_), .Y(_8597_) );
	AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_8597_), .B(_6879__bF_buf18), .Y(_6710__24_) );
	INVX1 INVX1_1481 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_25_), .Y(_8598_) );
	OAI21X1 OAI21X1_3630 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_8557__bF_buf2), .C(_6879__bF_buf17), .Y(_8599_) );
	AOI21X1 AOI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_8598_), .B(_8557__bF_buf1), .C(_8599_), .Y(_6710__25_) );
	OAI21X1 OAI21X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf11_bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_26_), .Y(_8600_) );
	OAI21X1 OAI21X1_3632 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_8557__bF_buf0), .C(_8600_), .Y(_8601_) );
	AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_8601_), .B(_6879__bF_buf16), .Y(_6710__26_) );
	INVX1 INVX1_1482 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_27_), .Y(_8602_) );
	OAI21X1 OAI21X1_3633 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_8557__bF_buf5), .C(_6879__bF_buf15), .Y(_8603_) );
	AOI21X1 AOI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_8602_), .B(_8557__bF_buf4), .C(_8603_), .Y(_6710__27_) );
	OAI21X1 OAI21X1_3634 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf10_bF_buf1), .B(_8554_), .C(csr_gpr_iu_csr_mideleg_28_), .Y(_8604_) );
	OAI21X1 OAI21X1_3635 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_8557__bF_buf3), .C(_8604_), .Y(_8605_) );
	AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_8605_), .B(_6879__bF_buf14), .Y(_6710__28_) );
	INVX1 INVX1_1483 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_29_), .Y(_8606_) );
	OAI21X1 OAI21X1_3636 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_8557__bF_buf2), .C(_6879__bF_buf13), .Y(_8607_) );
	AOI21X1 AOI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_8606_), .B(_8557__bF_buf1), .C(_8607_), .Y(_6710__29_) );
	NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_8556_), .Y(_8608_) );
	OAI21X1 OAI21X1_3637 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_30_), .B(_8556_), .C(_8608_), .Y(_8609_) );
	NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_8609_), .Y(_6710__30_) );
	INVX1 INVX1_1484 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_31_), .Y(_8610_) );
	OAI21X1 OAI21X1_3638 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf1), .B(_8557__bF_buf0), .C(_6879__bF_buf12), .Y(_8611_) );
	AOI21X1 AOI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_8610_), .B(_8557__bF_buf5), .C(_8611_), .Y(_6710__31_) );
	INVX1 INVX1_1485 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_0_), .Y(_8612_) );
	INVX1 INVX1_1486 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf2), .Y(_8613_) );
	NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_8613_), .Y(_8614_) );
	INVX4 INVX4_19 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .Y(_8615_) );
	NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_7424__bF_buf2), .Y(_8616_) );
	NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_8112_), .Y(_8617_) );
	INVX8 INVX8_77 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .Y(_8618_) );
	AOI22X1 AOI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(_7956_), .B(_8616__bF_buf8), .C(_7325_), .D(_8618__bF_buf6), .Y(_8619_) );
	OAI21X1 OAI21X1_3639 ( .gnd(gnd), .vdd(vdd), .A(_8616__bF_buf7), .B(_7303__bF_buf3_bF_buf1), .C(_6879__bF_buf11), .Y(_8620_) );
	AOI21X1 AOI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .B(_7303__bF_buf2), .C(_8620_), .Y(_8621_) );
	OAI22X1 OAI22X1_713 ( .gnd(gnd), .vdd(vdd), .A(_8612_), .B(_8621__bF_buf4), .C(rst_bF_buf67), .D(_8619_), .Y(_6722__0_) );
	INVX1 INVX1_1487 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_1_), .Y(_8622_) );
	AOI22X1 AOI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(_7964_), .B(_8616__bF_buf6), .C(_7329_), .D(_8618__bF_buf5), .Y(_8623_) );
	OAI22X1 OAI22X1_714 ( .gnd(gnd), .vdd(vdd), .A(_8622_), .B(_8621__bF_buf3), .C(rst_bF_buf66), .D(_8623_), .Y(_6722__1_) );
	INVX1 INVX1_1488 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_2_), .Y(_8624_) );
	AOI22X1 AOI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_8616__bF_buf5), .C(_7333_), .D(_8618__bF_buf4), .Y(_8625_) );
	OAI22X1 OAI22X1_715 ( .gnd(gnd), .vdd(vdd), .A(_8624_), .B(_8621__bF_buf2), .C(rst_bF_buf65), .D(_8625_), .Y(_6722__2_) );
	INVX1 INVX1_1489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_3_), .Y(_8626_) );
	AOI22X1 AOI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(_7970_), .B(_8616__bF_buf4), .C(_7336_), .D(_8618__bF_buf3), .Y(_8627_) );
	OAI22X1 OAI22X1_716 ( .gnd(gnd), .vdd(vdd), .A(_8626_), .B(_8621__bF_buf1), .C(rst_bF_buf64), .D(_8627_), .Y(_6722__3_) );
	INVX1 INVX1_1490 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_4_), .Y(_8628_) );
	AOI22X1 AOI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(_7973_), .B(_8616__bF_buf3), .C(_7339_), .D(_8618__bF_buf2), .Y(_8629_) );
	OAI22X1 OAI22X1_717 ( .gnd(gnd), .vdd(vdd), .A(_8628_), .B(_8621__bF_buf0), .C(rst_bF_buf63), .D(_8629_), .Y(_6722__4_) );
	INVX1 INVX1_1491 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_5_), .Y(_8630_) );
	AOI22X1 AOI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_8616__bF_buf2), .C(_7342_), .D(_8618__bF_buf1), .Y(_8631_) );
	OAI22X1 OAI22X1_718 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .B(_8621__bF_buf4), .C(rst_bF_buf62), .D(_8631_), .Y(_6722__5_) );
	INVX1 INVX1_1492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_6_), .Y(_8632_) );
	AOI22X1 AOI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_8616__bF_buf1), .C(_7345_), .D(_8618__bF_buf0), .Y(_8633_) );
	OAI22X1 OAI22X1_719 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .B(_8621__bF_buf3), .C(rst_bF_buf61), .D(_8633_), .Y(_6722__6_) );
	INVX1 INVX1_1493 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_7_), .Y(_8634_) );
	AOI22X1 AOI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(_7982_), .B(_8616__bF_buf0), .C(_7348_), .D(_8618__bF_buf6), .Y(_8635_) );
	OAI22X1 OAI22X1_720 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(_8621__bF_buf2), .C(rst_bF_buf60), .D(_8635_), .Y(_6722__7_) );
	INVX1 INVX1_1494 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_8_), .Y(_8636_) );
	AOI22X1 AOI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(_7985_), .B(_8616__bF_buf8), .C(_7351_), .D(_8618__bF_buf5), .Y(_8637_) );
	OAI22X1 OAI22X1_721 ( .gnd(gnd), .vdd(vdd), .A(_8636_), .B(_8621__bF_buf1), .C(rst_bF_buf59), .D(_8637_), .Y(_6722__8_) );
	INVX1 INVX1_1495 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_9_), .Y(_8638_) );
	AOI22X1 AOI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .B(_8616__bF_buf7), .C(_7354_), .D(_8618__bF_buf4), .Y(_8639_) );
	OAI22X1 OAI22X1_722 ( .gnd(gnd), .vdd(vdd), .A(_8638_), .B(_8621__bF_buf0), .C(rst_bF_buf58), .D(_8639_), .Y(_6722__9_) );
	INVX1 INVX1_1496 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_10_), .Y(_8640_) );
	AOI22X1 AOI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(_7991_), .B(_8616__bF_buf6), .C(_7357_), .D(_8618__bF_buf3), .Y(_8641_) );
	OAI22X1 OAI22X1_723 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8621__bF_buf4), .C(rst_bF_buf57), .D(_8641_), .Y(_6722__10_) );
	INVX1 INVX1_1497 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_11_), .Y(_8642_) );
	AOI22X1 AOI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(_7994_), .B(_8616__bF_buf5), .C(_7360_), .D(_8618__bF_buf2), .Y(_8643_) );
	OAI22X1 OAI22X1_724 ( .gnd(gnd), .vdd(vdd), .A(_8642_), .B(_8621__bF_buf3), .C(rst_bF_buf56), .D(_8643_), .Y(_6722__11_) );
	INVX1 INVX1_1498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_12_), .Y(_8644_) );
	AOI22X1 AOI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(_7997_), .B(_8616__bF_buf4), .C(_7363_), .D(_8618__bF_buf1), .Y(_8645_) );
	OAI22X1 OAI22X1_725 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .B(_8621__bF_buf2), .C(rst_bF_buf55), .D(_8645_), .Y(_6722__12_) );
	INVX1 INVX1_1499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_13_), .Y(_8646_) );
	AOI22X1 AOI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(_8000_), .B(_8616__bF_buf3), .C(_7492_), .D(_8618__bF_buf0), .Y(_8647_) );
	OAI22X1 OAI22X1_726 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_8621__bF_buf1), .C(rst_bF_buf54), .D(_8647_), .Y(_6722__13_) );
	INVX1 INVX1_1500 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_14_), .Y(_8648_) );
	AOI22X1 AOI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(_8003_), .B(_8616__bF_buf2), .C(_7370_), .D(_8618__bF_buf6), .Y(_8649_) );
	OAI22X1 OAI22X1_727 ( .gnd(gnd), .vdd(vdd), .A(_8648_), .B(_8621__bF_buf0), .C(rst_bF_buf53), .D(_8649_), .Y(_6722__14_) );
	INVX1 INVX1_1501 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_15_), .Y(_8650_) );
	AOI22X1 AOI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(_8006_), .B(_8616__bF_buf1), .C(_7501_), .D(_8618__bF_buf5), .Y(_8651_) );
	OAI22X1 OAI22X1_728 ( .gnd(gnd), .vdd(vdd), .A(_8650_), .B(_8621__bF_buf4), .C(rst_bF_buf52), .D(_8651_), .Y(_6722__15_) );
	INVX1 INVX1_1502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_16_), .Y(_8652_) );
	AOI22X1 AOI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(_8009_), .B(_8616__bF_buf0), .C(_7376_), .D(_8618__bF_buf4), .Y(_8653_) );
	OAI22X1 OAI22X1_729 ( .gnd(gnd), .vdd(vdd), .A(_8652_), .B(_8621__bF_buf3), .C(rst_bF_buf51), .D(_8653_), .Y(_6722__16_) );
	INVX1 INVX1_1503 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_17_), .Y(_8654_) );
	AOI22X1 AOI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_8616__bF_buf8), .C(_7510_), .D(_8618__bF_buf3), .Y(_8655_) );
	OAI22X1 OAI22X1_730 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_8621__bF_buf2), .C(rst_bF_buf50), .D(_8655_), .Y(_6722__17_) );
	INVX1 INVX1_1504 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_18_), .Y(_8656_) );
	AOI22X1 AOI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(_8015_), .B(_8616__bF_buf7), .C(_7382_), .D(_8618__bF_buf2), .Y(_8657_) );
	OAI22X1 OAI22X1_731 ( .gnd(gnd), .vdd(vdd), .A(_8656_), .B(_8621__bF_buf1), .C(rst_bF_buf49), .D(_8657_), .Y(_6722__18_) );
	INVX1 INVX1_1505 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_19_), .Y(_8658_) );
	AOI22X1 AOI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(_8018_), .B(_8616__bF_buf6), .C(_7519_), .D(_8618__bF_buf1), .Y(_8659_) );
	OAI22X1 OAI22X1_732 ( .gnd(gnd), .vdd(vdd), .A(_8658_), .B(_8621__bF_buf0), .C(rst_bF_buf48), .D(_8659_), .Y(_6722__19_) );
	INVX1 INVX1_1506 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_20_), .Y(_8660_) );
	AOI22X1 AOI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(_8021_), .B(_8616__bF_buf5), .C(_7388_), .D(_8618__bF_buf0), .Y(_8661_) );
	OAI22X1 OAI22X1_733 ( .gnd(gnd), .vdd(vdd), .A(_8660_), .B(_8621__bF_buf4), .C(rst_bF_buf47), .D(_8661_), .Y(_6722__20_) );
	INVX1 INVX1_1507 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_21_), .Y(_8662_) );
	AOI22X1 AOI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .B(_8616__bF_buf4), .C(_7528_), .D(_8618__bF_buf6), .Y(_8663_) );
	OAI22X1 OAI22X1_734 ( .gnd(gnd), .vdd(vdd), .A(_8662_), .B(_8621__bF_buf3), .C(rst_bF_buf46), .D(_8663_), .Y(_6722__21_) );
	INVX1 INVX1_1508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_22_), .Y(_8664_) );
	AOI22X1 AOI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(_8027_), .B(_8616__bF_buf3), .C(_7394_), .D(_8618__bF_buf5), .Y(_8665_) );
	OAI22X1 OAI22X1_735 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .B(_8621__bF_buf2), .C(rst_bF_buf45), .D(_8665_), .Y(_6722__22_) );
	INVX1 INVX1_1509 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_23_), .Y(_8666_) );
	AOI22X1 AOI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(_8616__bF_buf2), .C(_7537_), .D(_8618__bF_buf4), .Y(_8667_) );
	OAI22X1 OAI22X1_736 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8621__bF_buf1), .C(rst_bF_buf44), .D(_8667_), .Y(_6722__23_) );
	INVX1 INVX1_1510 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_24_), .Y(_8668_) );
	AOI22X1 AOI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(_8033_), .B(_8616__bF_buf1), .C(_7400_), .D(_8618__bF_buf3), .Y(_8669_) );
	OAI22X1 OAI22X1_737 ( .gnd(gnd), .vdd(vdd), .A(_8668_), .B(_8621__bF_buf0), .C(rst_bF_buf43), .D(_8669_), .Y(_6722__24_) );
	INVX1 INVX1_1511 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_25_), .Y(_8670_) );
	AOI22X1 AOI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8616__bF_buf0), .C(_7546_), .D(_8618__bF_buf2), .Y(_8671_) );
	OAI22X1 OAI22X1_738 ( .gnd(gnd), .vdd(vdd), .A(_8670_), .B(_8621__bF_buf4), .C(rst_bF_buf42), .D(_8671_), .Y(_6722__25_) );
	INVX1 INVX1_1512 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_26_), .Y(_8672_) );
	AOI22X1 AOI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(_8039_), .B(_8616__bF_buf8), .C(_7406_), .D(_8618__bF_buf1), .Y(_8673_) );
	OAI22X1 OAI22X1_739 ( .gnd(gnd), .vdd(vdd), .A(_8672_), .B(_8621__bF_buf3), .C(rst_bF_buf41), .D(_8673_), .Y(_6722__26_) );
	INVX1 INVX1_1513 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_27_), .Y(_8674_) );
	AOI22X1 AOI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(_8042_), .B(_8616__bF_buf7), .C(_7556_), .D(_8618__bF_buf0), .Y(_8675_) );
	OAI22X1 OAI22X1_740 ( .gnd(gnd), .vdd(vdd), .A(_8674_), .B(_8621__bF_buf2), .C(rst_bF_buf40), .D(_8675_), .Y(_6722__27_) );
	INVX1 INVX1_1514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_28_), .Y(_8676_) );
	AOI22X1 AOI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(_8045_), .B(_8616__bF_buf6), .C(_7412_), .D(_8618__bF_buf6), .Y(_8677_) );
	OAI22X1 OAI22X1_741 ( .gnd(gnd), .vdd(vdd), .A(_8676_), .B(_8621__bF_buf1), .C(rst_bF_buf39), .D(_8677_), .Y(_6722__28_) );
	INVX1 INVX1_1515 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_29_), .Y(_8678_) );
	AOI22X1 AOI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_8616__bF_buf5), .C(_7565_), .D(_8618__bF_buf5), .Y(_8679_) );
	OAI22X1 OAI22X1_742 ( .gnd(gnd), .vdd(vdd), .A(_8678_), .B(_8621__bF_buf0), .C(rst_bF_buf38), .D(_8679_), .Y(_6722__29_) );
	INVX1 INVX1_1516 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_30_), .Y(_8680_) );
	AOI22X1 AOI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_8616__bF_buf4), .C(_7417_), .D(_8618__bF_buf4), .Y(_8681_) );
	OAI22X1 OAI22X1_743 ( .gnd(gnd), .vdd(vdd), .A(_8680_), .B(_8621__bF_buf4), .C(rst_bF_buf37), .D(_8681_), .Y(_6722__30_) );
	INVX1 INVX1_1517 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_31_), .Y(_8682_) );
	AOI22X1 AOI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(_8054_), .B(_8616__bF_buf3), .C(_7574_), .D(_8618__bF_buf3), .Y(_8683_) );
	OAI22X1 OAI22X1_744 ( .gnd(gnd), .vdd(vdd), .A(_8682_), .B(_8621__bF_buf3), .C(rst_bF_buf36), .D(_8683_), .Y(_6722__31_) );
	NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_8161_), .Y(_8684_) );
	INVX1 INVX1_1518 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_0_), .Y(_8685_) );
	OAI21X1 OAI21X1_3640 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf3), .C(_8685_), .Y(_8686_) );
	OAI21X1 OAI21X1_3641 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_8684__bF_buf5), .C(_8686_), .Y(_8687_) );
	MUX2X1 MUX2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_8685_), .S(_8616__bF_buf2), .Y(_8688_) );
	OAI21X1 OAI21X1_3642 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf1), .B(_8688_), .C(_6879__bF_buf10), .Y(_8689_) );
	AOI21X1 AOI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_7303__bF_buf0), .C(_8689_), .Y(_6704__0_) );
	INVX1 INVX1_1519 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_1_), .Y(_8690_) );
	OAI21X1 OAI21X1_3643 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf2), .C(_8690_), .Y(_8691_) );
	OAI21X1 OAI21X1_3644 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_8684__bF_buf4), .C(_8691_), .Y(_8692_) );
	MUX2X1 MUX2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_7441_), .B(_8690_), .S(_8616__bF_buf1), .Y(_8693_) );
	OAI21X1 OAI21X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14_bF_buf0), .B(_8693_), .C(_6879__bF_buf9), .Y(_8694_) );
	AOI21X1 AOI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_8692_), .B(_7303__bF_buf13_bF_buf0), .C(_8694_), .Y(_6704__1_) );
	INVX1 INVX1_1520 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_2_), .Y(_8695_) );
	OAI21X1 OAI21X1_3646 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf4), .B(_7434__bF_buf1), .C(_8695_), .Y(_8696_) );
	OAI21X1 OAI21X1_3647 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_8684__bF_buf3), .C(_8696_), .Y(_8697_) );
	MUX2X1 MUX2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_8695_), .S(_8616__bF_buf0), .Y(_8698_) );
	OAI21X1 OAI21X1_3648 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12_bF_buf0), .B(_8698_), .C(_6879__bF_buf8), .Y(_8699_) );
	AOI21X1 AOI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .B(_7303__bF_buf11_bF_buf0), .C(_8699_), .Y(_6704__2_) );
	INVX1 INVX1_1521 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_3_), .Y(_8700_) );
	OAI21X1 OAI21X1_3649 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_7434__bF_buf0), .C(_8700_), .Y(_8701_) );
	OAI21X1 OAI21X1_3650 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_8684__bF_buf2), .C(_8701_), .Y(_8702_) );
	MUX2X1 MUX2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_8700_), .S(_8616__bF_buf8), .Y(_8703_) );
	OAI21X1 OAI21X1_3651 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf0), .B(_8703_), .C(_6879__bF_buf7), .Y(_8704_) );
	AOI21X1 AOI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_8702_), .B(_7303__bF_buf9_bF_buf0), .C(_8704_), .Y(_6704__3_) );
	INVX1 INVX1_1522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_4_), .Y(_8705_) );
	OAI21X1 OAI21X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf4), .C(_8705_), .Y(_8706_) );
	OAI21X1 OAI21X1_3653 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_8684__bF_buf1), .C(_8706_), .Y(_8707_) );
	MUX2X1 MUX2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_8705_), .S(_8616__bF_buf7), .Y(_8708_) );
	OAI21X1 OAI21X1_3654 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8_bF_buf0), .B(_8708_), .C(_6879__bF_buf6), .Y(_8709_) );
	AOI21X1 AOI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_8707_), .B(_7303__bF_buf7_bF_buf0), .C(_8709_), .Y(_6704__4_) );
	INVX1 INVX1_1523 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_5_), .Y(_8710_) );
	OAI21X1 OAI21X1_3655 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_7434__bF_buf3), .C(_8710_), .Y(_8711_) );
	OAI21X1 OAI21X1_3656 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_8684__bF_buf0), .C(_8711_), .Y(_8712_) );
	MUX2X1 MUX2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .B(_8710_), .S(_8616__bF_buf6), .Y(_8713_) );
	OAI21X1 OAI21X1_3657 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6_bF_buf0), .B(_8713_), .C(_6879__bF_buf5), .Y(_8714_) );
	AOI21X1 AOI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_8712_), .B(_7303__bF_buf5_bF_buf0), .C(_8714_), .Y(_6704__5_) );
	INVX1 INVX1_1524 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_6_), .Y(_8715_) );
	OAI21X1 OAI21X1_3658 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf2), .C(_8715_), .Y(_8716_) );
	OAI21X1 OAI21X1_3659 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_8684__bF_buf5), .C(_8716_), .Y(_8717_) );
	MUX2X1 MUX2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_8715_), .S(_8616__bF_buf5), .Y(_8718_) );
	OAI21X1 OAI21X1_3660 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4_bF_buf0), .B(_8718_), .C(_6879__bF_buf4), .Y(_8719_) );
	AOI21X1 AOI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_8717_), .B(_7303__bF_buf3_bF_buf0), .C(_8719_), .Y(_6704__6_) );
	INVX1 INVX1_1525 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_7_), .Y(_8720_) );
	OAI21X1 OAI21X1_3661 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf1), .C(_8720_), .Y(_8721_) );
	OAI21X1 OAI21X1_3662 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_8684__bF_buf4), .C(_8721_), .Y(_8722_) );
	MUX2X1 MUX2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .B(_8720_), .S(_8616__bF_buf4), .Y(_8723_) );
	OAI21X1 OAI21X1_3663 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf2), .B(_8723_), .C(_6879__bF_buf3), .Y(_8724_) );
	AOI21X1 AOI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_8722_), .B(_7303__bF_buf1), .C(_8724_), .Y(_6704__7_) );
	INVX1 INVX1_1526 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_8_), .Y(_8725_) );
	OAI21X1 OAI21X1_3664 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf4), .B(_7434__bF_buf0), .C(_8725_), .Y(_8726_) );
	OAI21X1 OAI21X1_3665 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_8684__bF_buf3), .C(_8726_), .Y(_8727_) );
	MUX2X1 MUX2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_7469_), .B(_8725_), .S(_8616__bF_buf3), .Y(_8728_) );
	OAI21X1 OAI21X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf0), .B(_8728_), .C(_6879__bF_buf2), .Y(_8729_) );
	AOI21X1 AOI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_8727_), .B(_7303__bF_buf14_bF_buf3), .C(_8729_), .Y(_6704__8_) );
	INVX1 INVX1_1527 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_9_), .Y(_8730_) );
	OAI21X1 OAI21X1_3667 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_7434__bF_buf4), .C(_8730_), .Y(_8731_) );
	OAI21X1 OAI21X1_3668 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_8684__bF_buf2), .C(_8731_), .Y(_8732_) );
	MUX2X1 MUX2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_8730_), .S(_8616__bF_buf2), .Y(_8733_) );
	OAI21X1 OAI21X1_3669 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13_bF_buf3), .B(_8733_), .C(_6879__bF_buf1), .Y(_8734_) );
	AOI21X1 AOI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .B(_7303__bF_buf12_bF_buf3), .C(_8734_), .Y(_6704__9_) );
	INVX1 INVX1_1528 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_10_), .Y(_8735_) );
	OAI21X1 OAI21X1_3670 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf3), .C(_8735_), .Y(_8736_) );
	OAI21X1 OAI21X1_3671 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_8684__bF_buf1), .C(_8736_), .Y(_8737_) );
	MUX2X1 MUX2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_7477_), .B(_8735_), .S(_8616__bF_buf1), .Y(_8738_) );
	OAI21X1 OAI21X1_3672 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11_bF_buf3), .B(_8738_), .C(_6879__bF_buf0), .Y(_8739_) );
	AOI21X1 AOI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_8737_), .B(_7303__bF_buf10_bF_buf3), .C(_8739_), .Y(_6704__10_) );
	INVX1 INVX1_1529 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_11_), .Y(_8740_) );
	OAI21X1 OAI21X1_3673 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_7434__bF_buf2), .C(_8740_), .Y(_8741_) );
	OAI21X1 OAI21X1_3674 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .B(_8684__bF_buf0), .C(_8741_), .Y(_8742_) );
	MUX2X1 MUX2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .B(_8740_), .S(_8616__bF_buf0), .Y(_8743_) );
	OAI21X1 OAI21X1_3675 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9_bF_buf3), .B(_8743_), .C(_6879__bF_buf42), .Y(_8744_) );
	AOI21X1 AOI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_7303__bF_buf8_bF_buf3), .C(_8744_), .Y(_6704__11_) );
	INVX1 INVX1_1530 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_12_), .Y(_8745_) );
	OAI21X1 OAI21X1_3676 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf1), .C(_8745_), .Y(_8746_) );
	OAI21X1 OAI21X1_3677 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_8684__bF_buf5), .C(_8746_), .Y(_8747_) );
	MUX2X1 MUX2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_8745_), .S(_8616__bF_buf8), .Y(_8748_) );
	OAI21X1 OAI21X1_3678 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7_bF_buf3), .B(_8748_), .C(_6879__bF_buf41), .Y(_8749_) );
	AOI21X1 AOI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_7303__bF_buf6_bF_buf3), .C(_8749_), .Y(_6704__12_) );
	INVX1 INVX1_1531 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_13_), .Y(_8750_) );
	OAI21X1 OAI21X1_3679 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf0), .C(_8750_), .Y(_8751_) );
	OAI21X1 OAI21X1_3680 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_8684__bF_buf4), .C(_8751_), .Y(_8752_) );
	MUX2X1 MUX2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_8750_), .S(_8616__bF_buf7), .Y(_8753_) );
	OAI21X1 OAI21X1_3681 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5_bF_buf3), .B(_8753_), .C(_6879__bF_buf40), .Y(_8754_) );
	AOI21X1 AOI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_8752_), .B(_7303__bF_buf4_bF_buf3), .C(_8754_), .Y(_6704__13_) );
	INVX1 INVX1_1532 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_14_), .Y(_8755_) );
	OAI21X1 OAI21X1_3682 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf4), .B(_7434__bF_buf4), .C(_8755_), .Y(_8756_) );
	OAI21X1 OAI21X1_3683 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_8684__bF_buf3), .C(_8756_), .Y(_8757_) );
	MUX2X1 MUX2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_7495_), .B(_8755_), .S(_8616__bF_buf6), .Y(_8758_) );
	OAI21X1 OAI21X1_3684 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3_bF_buf3), .B(_8758_), .C(_6879__bF_buf39), .Y(_8759_) );
	AOI21X1 AOI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_7303__bF_buf2), .C(_8759_), .Y(_6704__14_) );
	INVX1 INVX1_1533 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_15_), .Y(_8760_) );
	OAI21X1 OAI21X1_3685 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_7434__bF_buf3), .C(_8760_), .Y(_8761_) );
	OAI21X1 OAI21X1_3686 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf0), .B(_8684__bF_buf2), .C(_8761_), .Y(_8762_) );
	MUX2X1 MUX2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_8760_), .S(_8616__bF_buf5), .Y(_8763_) );
	OAI21X1 OAI21X1_3687 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf1), .B(_8763_), .C(_6879__bF_buf38), .Y(_8764_) );
	AOI21X1 AOI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_8762_), .B(_7303__bF_buf0), .C(_8764_), .Y(_6704__15_) );
	INVX1 INVX1_1534 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_16_), .Y(_8765_) );
	OAI21X1 OAI21X1_3688 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf2), .C(_8765_), .Y(_8766_) );
	OAI21X1 OAI21X1_3689 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_8684__bF_buf1), .C(_8766_), .Y(_8767_) );
	MUX2X1 MUX2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .B(_8765_), .S(_8616__bF_buf4), .Y(_8768_) );
	OAI21X1 OAI21X1_3690 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14_bF_buf2), .B(_8768_), .C(_6879__bF_buf37), .Y(_8769_) );
	AOI21X1 AOI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_8767_), .B(_7303__bF_buf13_bF_buf2), .C(_8769_), .Y(_6704__16_) );
	INVX1 INVX1_1535 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_17_), .Y(_8770_) );
	OAI21X1 OAI21X1_3691 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_7434__bF_buf1), .C(_8770_), .Y(_8771_) );
	OAI21X1 OAI21X1_3692 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf1), .B(_8684__bF_buf0), .C(_8771_), .Y(_8772_) );
	MUX2X1 MUX2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_8770_), .S(_8616__bF_buf3), .Y(_8773_) );
	OAI21X1 OAI21X1_3693 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12_bF_buf2), .B(_8773_), .C(_6879__bF_buf36), .Y(_8774_) );
	AOI21X1 AOI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .B(_7303__bF_buf11_bF_buf2), .C(_8774_), .Y(_6704__17_) );
	INVX1 INVX1_1536 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_18_), .Y(_8775_) );
	OAI21X1 OAI21X1_3694 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf0), .C(_8775_), .Y(_8776_) );
	OAI21X1 OAI21X1_3695 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_8684__bF_buf5), .C(_8776_), .Y(_8777_) );
	MUX2X1 MUX2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_7513_), .B(_8775_), .S(_8616__bF_buf2), .Y(_8778_) );
	OAI21X1 OAI21X1_3696 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf2), .B(_8778_), .C(_6879__bF_buf35), .Y(_8779_) );
	AOI21X1 AOI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .B(_7303__bF_buf9_bF_buf2), .C(_8779_), .Y(_6704__18_) );
	INVX1 INVX1_1537 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_19_), .Y(_8780_) );
	OAI21X1 OAI21X1_3697 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf4), .C(_8780_), .Y(_8781_) );
	OAI21X1 OAI21X1_3698 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf2), .B(_8684__bF_buf4), .C(_8781_), .Y(_8782_) );
	MUX2X1 MUX2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_7517_), .B(_8780_), .S(_8616__bF_buf1), .Y(_8783_) );
	OAI21X1 OAI21X1_3699 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8_bF_buf2), .B(_8783_), .C(_6879__bF_buf34), .Y(_8784_) );
	AOI21X1 AOI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .B(_7303__bF_buf7_bF_buf2), .C(_8784_), .Y(_6704__19_) );
	INVX1 INVX1_1538 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_20_), .Y(_8785_) );
	OAI21X1 OAI21X1_3700 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf4), .B(_7434__bF_buf3), .C(_8785_), .Y(_8786_) );
	OAI21X1 OAI21X1_3701 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_8684__bF_buf3), .C(_8786_), .Y(_8787_) );
	MUX2X1 MUX2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_7522_), .B(_8785_), .S(_8616__bF_buf0), .Y(_8788_) );
	OAI21X1 OAI21X1_3702 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6_bF_buf2), .B(_8788_), .C(_6879__bF_buf33), .Y(_8789_) );
	AOI21X1 AOI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_8787_), .B(_7303__bF_buf5_bF_buf2), .C(_8789_), .Y(_6704__20_) );
	INVX1 INVX1_1539 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_21_), .Y(_8790_) );
	OAI21X1 OAI21X1_3703 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_7434__bF_buf2), .C(_8790_), .Y(_8791_) );
	OAI21X1 OAI21X1_3704 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf2), .B(_8684__bF_buf2), .C(_8791_), .Y(_8792_) );
	MUX2X1 MUX2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_7526_), .B(_8790_), .S(_8616__bF_buf8), .Y(_8793_) );
	OAI21X1 OAI21X1_3705 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf4_bF_buf2), .B(_8793_), .C(_6879__bF_buf32), .Y(_8794_) );
	AOI21X1 AOI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .B(_7303__bF_buf3_bF_buf2), .C(_8794_), .Y(_6704__21_) );
	INVX1 INVX1_1540 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_22_), .Y(_8795_) );
	OAI21X1 OAI21X1_3706 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf1), .C(_8795_), .Y(_8796_) );
	OAI21X1 OAI21X1_3707 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_8684__bF_buf1), .C(_8796_), .Y(_8797_) );
	MUX2X1 MUX2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_7531_), .B(_8795_), .S(_8616__bF_buf7), .Y(_8798_) );
	OAI21X1 OAI21X1_3708 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf2), .B(_8798_), .C(_6879__bF_buf31), .Y(_8799_) );
	AOI21X1 AOI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_7303__bF_buf1), .C(_8799_), .Y(_6704__22_) );
	INVX1 INVX1_1541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_23_), .Y(_8800_) );
	OAI21X1 OAI21X1_3709 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_7434__bF_buf0), .C(_8800_), .Y(_8801_) );
	OAI21X1 OAI21X1_3710 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf0), .B(_8684__bF_buf0), .C(_8801_), .Y(_8802_) );
	MUX2X1 MUX2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_7535_), .B(_8800_), .S(_8616__bF_buf6), .Y(_8803_) );
	OAI21X1 OAI21X1_3711 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf0), .B(_8803_), .C(_6879__bF_buf30), .Y(_8804_) );
	AOI21X1 AOI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_7303__bF_buf14_bF_buf1), .C(_8804_), .Y(_6704__23_) );
	INVX1 INVX1_1542 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_24_), .Y(_8805_) );
	OAI21X1 OAI21X1_3712 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf4), .C(_8805_), .Y(_8806_) );
	OAI21X1 OAI21X1_3713 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_8684__bF_buf5), .C(_8806_), .Y(_8807_) );
	MUX2X1 MUX2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .B(_8805_), .S(_8616__bF_buf5), .Y(_8808_) );
	OAI21X1 OAI21X1_3714 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf13_bF_buf1), .B(_8808_), .C(_6879__bF_buf29), .Y(_8809_) );
	AOI21X1 AOI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_8807_), .B(_7303__bF_buf12_bF_buf1), .C(_8809_), .Y(_6704__24_) );
	INVX1 INVX1_1543 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_25_), .Y(_8810_) );
	OAI21X1 OAI21X1_3715 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf3), .C(_8810_), .Y(_8811_) );
	OAI21X1 OAI21X1_3716 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf2), .B(_8684__bF_buf4), .C(_8811_), .Y(_8812_) );
	MUX2X1 MUX2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_7544_), .B(_8810_), .S(_8616__bF_buf4), .Y(_8813_) );
	OAI21X1 OAI21X1_3717 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11_bF_buf1), .B(_8813_), .C(_6879__bF_buf28), .Y(_8814_) );
	AOI21X1 AOI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_7303__bF_buf10_bF_buf1), .C(_8814_), .Y(_6704__25_) );
	INVX1 INVX1_1544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_26_), .Y(_8815_) );
	OAI21X1 OAI21X1_3718 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf4), .B(_7434__bF_buf2), .C(_8815_), .Y(_8816_) );
	OAI21X1 OAI21X1_3719 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .B(_8684__bF_buf3), .C(_8816_), .Y(_8817_) );
	MUX2X1 MUX2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_7549_), .B(_8815_), .S(_8616__bF_buf3), .Y(_8818_) );
	OAI21X1 OAI21X1_3720 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9_bF_buf1), .B(_8818_), .C(_6879__bF_buf27), .Y(_8819_) );
	AOI21X1 AOI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_7303__bF_buf8_bF_buf1), .C(_8819_), .Y(_6704__26_) );
	INVX1 INVX1_1545 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_27_), .Y(_8820_) );
	OAI21X1 OAI21X1_3721 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf3), .B(_7434__bF_buf1), .C(_8820_), .Y(_8821_) );
	OAI21X1 OAI21X1_3722 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf2), .B(_8684__bF_buf2), .C(_8821_), .Y(_8822_) );
	MUX2X1 MUX2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_7553_), .B(_8820_), .S(_8616__bF_buf2), .Y(_8823_) );
	OAI21X1 OAI21X1_3723 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7_bF_buf1), .B(_8823_), .C(_6879__bF_buf26), .Y(_8824_) );
	AOI21X1 AOI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_8822_), .B(_7303__bF_buf6_bF_buf1), .C(_8824_), .Y(_6704__27_) );
	INVX1 INVX1_1546 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_28_), .Y(_8825_) );
	OAI21X1 OAI21X1_3724 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf0), .C(_8825_), .Y(_8826_) );
	OAI21X1 OAI21X1_3725 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_8684__bF_buf1), .C(_8826_), .Y(_8827_) );
	MUX2X1 MUX2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_7559_), .B(_8825_), .S(_8616__bF_buf1), .Y(_8828_) );
	OAI21X1 OAI21X1_3726 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5_bF_buf1), .B(_8828_), .C(_6879__bF_buf25), .Y(_8829_) );
	AOI21X1 AOI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_8827_), .B(_7303__bF_buf4_bF_buf1), .C(_8829_), .Y(_6704__28_) );
	INVX1 INVX1_1547 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_29_), .Y(_8830_) );
	OAI21X1 OAI21X1_3727 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_7434__bF_buf4), .C(_8830_), .Y(_8831_) );
	OAI21X1 OAI21X1_3728 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf2), .B(_8684__bF_buf0), .C(_8831_), .Y(_8832_) );
	MUX2X1 MUX2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .B(_8830_), .S(_8616__bF_buf0), .Y(_8833_) );
	OAI21X1 OAI21X1_3729 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3_bF_buf1), .B(_8833_), .C(_6879__bF_buf24), .Y(_8834_) );
	AOI21X1 AOI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_8832_), .B(_7303__bF_buf2), .C(_8834_), .Y(_6704__29_) );
	INVX1 INVX1_1548 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_30_), .Y(_8835_) );
	OAI21X1 OAI21X1_3730 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf0), .B(_7434__bF_buf3), .C(_8835_), .Y(_8836_) );
	OAI21X1 OAI21X1_3731 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_8684__bF_buf5), .C(_8836_), .Y(_8837_) );
	MUX2X1 MUX2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_7568_), .B(_8835_), .S(_8616__bF_buf8), .Y(_8838_) );
	OAI21X1 OAI21X1_3732 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf1), .B(_8838_), .C(_6879__bF_buf23), .Y(_8839_) );
	AOI21X1 AOI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_8837_), .B(_7303__bF_buf0), .C(_8839_), .Y(_6704__30_) );
	INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_31_), .Y(_8840_) );
	OAI21X1 OAI21X1_3733 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf5), .B(_7434__bF_buf2), .C(_8840_), .Y(_8841_) );
	OAI21X1 OAI21X1_3734 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf0), .B(_8684__bF_buf4), .C(_8841_), .Y(_8842_) );
	MUX2X1 MUX2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_7572_), .B(_8840_), .S(_8616__bF_buf7), .Y(_8843_) );
	OAI21X1 OAI21X1_3735 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14_bF_buf0), .B(_8843_), .C(_6879__bF_buf22), .Y(_8844_) );
	AOI21X1 AOI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_8842_), .B(_7303__bF_buf13_bF_buf0), .C(_8844_), .Y(_6704__31_) );
	INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .Y(_8845_) );
	NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_8230_), .Y(_8846_) );
	INVX8 INVX8_78 ( .gnd(gnd), .vdd(vdd), .A(_8846__bF_buf3), .Y(_8847_) );
	INVX1 INVX1_1549 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_0_), .Y(_8848_) );
	OAI21X1 OAI21X1_3736 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_8230_), .C(_8848_), .Y(_8849_) );
	OAI21X1 OAI21X1_3737 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_8847__bF_buf7), .C(_8849_), .Y(_8850_) );
	MUX2X1 MUX2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_8848_), .S(_8616__bF_buf6), .Y(_8851_) );
	OAI21X1 OAI21X1_3738 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12_bF_buf0), .B(_8851_), .C(_6879__bF_buf21), .Y(_8852_) );
	AOI21X1 AOI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_8850_), .B(_7303__bF_buf11_bF_buf0), .C(_8852_), .Y(_6709__0_) );
	INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_1_), .Y(_8853_) );
	OAI21X1 OAI21X1_3739 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_8230_), .C(_8853_), .Y(_8854_) );
	OAI21X1 OAI21X1_3740 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_8847__bF_buf6), .C(_8854_), .Y(_8855_) );
	MUX2X1 MUX2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_8853_), .S(_8616__bF_buf5), .Y(_8856_) );
	OAI21X1 OAI21X1_3741 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf0), .B(_8856_), .C(_6879__bF_buf20), .Y(_8857_) );
	AOI21X1 AOI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_7303__bF_buf9_bF_buf0), .C(_8857_), .Y(_6709__1_) );
	INVX1 INVX1_1550 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_2_), .Y(_8858_) );
	AOI21X1 AOI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf5), .B(_8858_), .C(_7304__bF_buf9_bF_buf1), .Y(_8859_) );
	OAI21X1 OAI21X1_3742 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_8847__bF_buf4), .C(_8859_), .Y(_8860_) );
	INVX8 INVX8_79 ( .gnd(gnd), .vdd(vdd), .A(_8616__bF_buf4), .Y(_8861_) );
	AOI21X1 AOI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_8858_), .C(_7303__bF_buf8_bF_buf0), .Y(_8862_) );
	OAI21X1 OAI21X1_3743 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_7621_), .C(_8862_), .Y(_8863_) );
	AOI21X1 AOI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8860_), .C(rst_bF_buf35), .Y(_6709__2_) );
	INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_3_), .Y(_8864_) );
	AOI21X1 AOI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf3), .B(_8864_), .C(_7304__bF_buf8_bF_buf1), .Y(_8865_) );
	OAI21X1 OAI21X1_3744 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_8847__bF_buf2), .C(_8865_), .Y(_8866_) );
	AOI21X1 AOI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_8864_), .C(_7303__bF_buf7_bF_buf0), .Y(_8867_) );
	OAI21X1 OAI21X1_3745 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_7637_), .C(_8867_), .Y(_8868_) );
	AOI21X1 AOI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .B(_8866_), .C(rst_bF_buf34), .Y(_6709__3_) );
	INVX1 INVX1_1551 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_4_), .Y(_8869_) );
	AOI21X1 AOI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf1), .B(_8869_), .C(_7304__bF_buf7_bF_buf1), .Y(_8870_) );
	OAI21X1 OAI21X1_3746 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_8847__bF_buf0), .C(_8870_), .Y(_8871_) );
	AOI21X1 AOI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_8869_), .C(_7303__bF_buf6_bF_buf0), .Y(_8872_) );
	OAI21X1 OAI21X1_3747 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_7647_), .C(_8872_), .Y(_8873_) );
	AOI21X1 AOI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .B(_8871_), .C(rst_bF_buf33), .Y(_6709__4_) );
	INVX1 INVX1_1552 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_5_), .Y(_8874_) );
	AOI21X1 AOI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf7), .B(_8874_), .C(_7304__bF_buf6_bF_buf1), .Y(_8875_) );
	OAI21X1 OAI21X1_3748 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_8847__bF_buf6), .C(_8875_), .Y(_8876_) );
	AOI21X1 AOI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_8874_), .C(_7303__bF_buf5_bF_buf0), .Y(_8877_) );
	OAI21X1 OAI21X1_3749 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_7658_), .C(_8877_), .Y(_8878_) );
	AOI21X1 AOI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_8878_), .B(_8876_), .C(rst_bF_buf32), .Y(_6709__5_) );
	OAI21X1 OAI21X1_3750 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_7424__bF_buf1), .C(csr_gpr_iu_csr_mepc_6_), .Y(_8879_) );
	OAI21X1 OAI21X1_3751 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_7667_), .C(_8879_), .Y(_8880_) );
	OAI21X1 OAI21X1_3752 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf2), .C(_8880_), .Y(_8881_) );
	INVX1 INVX1_1553 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_6_), .Y(_8882_) );
	AOI21X1 AOI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf5), .B(_8882_), .C(_7304__bF_buf5), .Y(_8883_) );
	OAI21X1 OAI21X1_3753 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_8847__bF_buf4), .C(_8883_), .Y(_8884_) );
	AOI21X1 AOI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_8884_), .C(rst_bF_buf31), .Y(_6709__6_) );
	INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_7_), .Y(_8885_) );
	AOI21X1 AOI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_8885_), .C(_7303__bF_buf4_bF_buf0), .Y(_8886_) );
	OAI21X1 OAI21X1_3754 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_7677_), .C(_8886_), .Y(_8887_) );
	AOI21X1 AOI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf3), .B(_8885_), .C(_7304__bF_buf4), .Y(_8888_) );
	OAI21X1 OAI21X1_3755 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_8847__bF_buf2), .C(_8888_), .Y(_8889_) );
	AOI21X1 AOI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_8887_), .B(_8889_), .C(rst_bF_buf30), .Y(_6709__7_) );
	INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_8_), .Y(_8890_) );
	OAI21X1 OAI21X1_3756 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_7424__bF_buf0), .C(_8890_), .Y(_8891_) );
	OAI21X1 OAI21X1_3757 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_7690_), .C(_8891_), .Y(_8892_) );
	NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_7583__bF_buf3), .B(_8111__bF_buf4), .Y(_8893_) );
	NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_8890_), .B(_8893_), .Y(_8894_) );
	OAI21X1 OAI21X1_3758 ( .gnd(gnd), .vdd(vdd), .A(_6927_), .B(_8847__bF_buf1), .C(_7303__bF_buf3_bF_buf0), .Y(_8895_) );
	OAI21X1 OAI21X1_3759 ( .gnd(gnd), .vdd(vdd), .A(_8894_), .B(_8895_), .C(_6879__bF_buf19), .Y(_8896_) );
	AOI21X1 AOI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_8892_), .B(_7304__bF_buf3), .C(_8896_), .Y(_6709__8_) );
	INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_9_), .Y(_8897_) );
	AOI21X1 AOI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf0), .B(_8897_), .C(_7304__bF_buf2), .Y(_8898_) );
	OAI21X1 OAI21X1_3760 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_8847__bF_buf7), .C(_8898_), .Y(_8899_) );
	AOI21X1 AOI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_8897_), .C(_7303__bF_buf2), .Y(_8900_) );
	OAI21X1 OAI21X1_3761 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_7701_), .C(_8900_), .Y(_8901_) );
	AOI21X1 AOI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_8901_), .B(_8899_), .C(rst_bF_buf29), .Y(_6709__9_) );
	INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_10_), .Y(_8902_) );
	AOI21X1 AOI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf6), .B(_8902_), .C(_7304__bF_buf1), .Y(_8903_) );
	OAI21X1 OAI21X1_3762 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_8847__bF_buf5), .C(_8903_), .Y(_8904_) );
	AOI21X1 AOI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_8902_), .C(_7303__bF_buf1), .Y(_8905_) );
	OAI21X1 OAI21X1_3763 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_7715_), .C(_8905_), .Y(_8906_) );
	AOI21X1 AOI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_8906_), .B(_8904_), .C(rst_bF_buf28), .Y(_6709__10_) );
	INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_11_), .Y(_8907_) );
	AOI21X1 AOI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_8907_), .C(_7303__bF_buf0), .Y(_8908_) );
	OAI21X1 OAI21X1_3764 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_7727_), .C(_8908_), .Y(_8909_) );
	AOI21X1 AOI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf4), .B(_8907_), .C(_7304__bF_buf0), .Y(_8910_) );
	OAI21X1 OAI21X1_3765 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .B(_8847__bF_buf3), .C(_8910_), .Y(_8911_) );
	AOI21X1 AOI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_8911_), .C(rst_bF_buf27), .Y(_6709__11_) );
	INVX1 INVX1_1554 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_12_), .Y(_8912_) );
	OAI21X1 OAI21X1_3766 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_7424__bF_buf3), .C(_8912_), .Y(_8913_) );
	OAI21X1 OAI21X1_3767 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_7734_), .C(_8913_), .Y(_8914_) );
	NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_8912_), .B(_8893_), .Y(_8915_) );
	OAI21X1 OAI21X1_3768 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_8847__bF_buf2), .C(_7303__bF_buf14_bF_buf3), .Y(_8916_) );
	OAI21X1 OAI21X1_3769 ( .gnd(gnd), .vdd(vdd), .A(_8915_), .B(_8916_), .C(_6879__bF_buf18), .Y(_8917_) );
	AOI21X1 AOI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_8914_), .B(_7304__bF_buf14_bF_buf0), .C(_8917_), .Y(_6709__12_) );
	INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_13_), .Y(_8918_) );
	AOI21X1 AOI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf1), .B(_8918_), .C(_7304__bF_buf13_bF_buf0), .Y(_8919_) );
	OAI21X1 OAI21X1_3770 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf2), .B(_8847__bF_buf0), .C(_8919_), .Y(_8920_) );
	OAI21X1 OAI21X1_3771 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_7744_), .C(_8616__bF_buf3), .Y(_8921_) );
	AOI21X1 AOI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_8918_), .C(_7303__bF_buf13_bF_buf3), .Y(_8922_) );
	NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_8922_), .B(_8921_), .Y(_8923_) );
	AOI21X1 AOI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_8920_), .C(rst_bF_buf26), .Y(_6709__13_) );
	OAI21X1 OAI21X1_3772 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .B(_7757_), .C(_8616__bF_buf2), .Y(_8924_) );
	OAI21X1 OAI21X1_3773 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_14_), .B(_8616__bF_buf1), .C(_8924_), .Y(_8925_) );
	NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_8847__bF_buf7), .Y(_8926_) );
	INVX1 INVX1_1555 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_14_), .Y(_8927_) );
	OAI21X1 OAI21X1_3774 ( .gnd(gnd), .vdd(vdd), .A(_8927_), .B(_8893_), .C(_7303__bF_buf12_bF_buf3), .Y(_8928_) );
	OAI21X1 OAI21X1_3775 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(_8926_), .C(_6879__bF_buf17), .Y(_8929_) );
	AOI21X1 AOI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_8925_), .B(_7304__bF_buf12_bF_buf0), .C(_8929_), .Y(_6709__14_) );
	INVX1 INVX1_1556 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_15_), .Y(_8930_) );
	AOI21X1 AOI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf6), .B(_8930_), .C(_7304__bF_buf11_bF_buf0), .Y(_8931_) );
	OAI21X1 OAI21X1_3776 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf3), .B(_8847__bF_buf5), .C(_8931_), .Y(_8932_) );
	AOI21X1 AOI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_8930_), .C(_7303__bF_buf11_bF_buf3), .Y(_8933_) );
	OAI21X1 OAI21X1_3777 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_7767_), .C(_8933_), .Y(_8934_) );
	AOI21X1 AOI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_8934_), .B(_8932_), .C(rst_bF_buf25), .Y(_6709__15_) );
	INVX1 INVX1_1557 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_16_), .Y(_8935_) );
	AOI21X1 AOI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf4), .B(_8935_), .C(_7304__bF_buf10_bF_buf0), .Y(_8936_) );
	OAI21X1 OAI21X1_3778 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_8847__bF_buf3), .C(_8936_), .Y(_8937_) );
	OAI21X1 OAI21X1_3779 ( .gnd(gnd), .vdd(vdd), .A(_7778_), .B(_7774_), .C(_8616__bF_buf0), .Y(_8938_) );
	AOI21X1 AOI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_8935_), .C(_7303__bF_buf10_bF_buf3), .Y(_8939_) );
	NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_8939_), .B(_8938_), .Y(_8940_) );
	AOI21X1 AOI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(_8937_), .C(rst_bF_buf24), .Y(_6709__16_) );
	INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_17_), .Y(_8941_) );
	AOI21X1 AOI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf2), .B(_8941_), .C(_7304__bF_buf9_bF_buf0), .Y(_8942_) );
	OAI21X1 OAI21X1_3780 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf0), .B(_8847__bF_buf1), .C(_8942_), .Y(_8943_) );
	OAI21X1 OAI21X1_3781 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_7786_), .C(_8616__bF_buf8), .Y(_8944_) );
	AOI21X1 AOI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_8941_), .C(_7303__bF_buf9_bF_buf3), .Y(_8945_) );
	NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_8945_), .B(_8944_), .Y(_8946_) );
	AOI21X1 AOI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_8946_), .B(_8943_), .C(rst_bF_buf23), .Y(_6709__17_) );
	INVX1 INVX1_1558 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_18_), .Y(_8947_) );
	AOI21X1 AOI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf0), .B(_8947_), .C(_7304__bF_buf8_bF_buf0), .Y(_8948_) );
	OAI21X1 OAI21X1_3782 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_8847__bF_buf7), .C(_8948_), .Y(_8949_) );
	AOI21X1 AOI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_8947_), .C(_7303__bF_buf8_bF_buf3), .Y(_8950_) );
	OAI21X1 OAI21X1_3783 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_7801_), .C(_8950_), .Y(_8951_) );
	AOI21X1 AOI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(_8949_), .C(rst_bF_buf22), .Y(_6709__18_) );
	INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_19_), .Y(_8952_) );
	AOI21X1 AOI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf6), .B(_8952_), .C(_7304__bF_buf7_bF_buf0), .Y(_8953_) );
	OAI21X1 OAI21X1_3784 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf1), .B(_8847__bF_buf5), .C(_8953_), .Y(_8954_) );
	AOI21X1 AOI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_8952_), .C(_7303__bF_buf7_bF_buf3), .Y(_8955_) );
	OAI21X1 OAI21X1_3785 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_7812_), .C(_8955_), .Y(_8956_) );
	AOI21X1 AOI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_8956_), .B(_8954_), .C(rst_bF_buf21), .Y(_6709__19_) );
	INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_20_), .Y(_8957_) );
	AOI21X1 AOI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf4), .B(_8957_), .C(_7304__bF_buf6_bF_buf0), .Y(_8958_) );
	OAI21X1 OAI21X1_3786 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_8847__bF_buf3), .C(_8958_), .Y(_8959_) );
	AOI21X1 AOI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_8957_), .C(_7303__bF_buf6_bF_buf3), .Y(_8960_) );
	OAI21X1 OAI21X1_3787 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_7821_), .C(_8960_), .Y(_8961_) );
	AOI21X1 AOI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_8961_), .B(_8959_), .C(rst_bF_buf20), .Y(_6709__20_) );
	INVX1 INVX1_1559 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_21_), .Y(_8962_) );
	AOI21X1 AOI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf2), .B(_8962_), .C(_7304__bF_buf5), .Y(_8963_) );
	OAI21X1 OAI21X1_3788 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf1), .B(_8847__bF_buf1), .C(_8963_), .Y(_8964_) );
	AOI21X1 AOI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_8962_), .C(_7303__bF_buf5_bF_buf3), .Y(_8965_) );
	OAI21X1 OAI21X1_3789 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_7831_), .C(_8965_), .Y(_8966_) );
	AOI21X1 AOI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(_8964_), .C(rst_bF_buf19), .Y(_6709__21_) );
	INVX1 INVX1_1560 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_22_), .Y(_8967_) );
	AOI21X1 AOI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf0), .B(_8967_), .C(_7304__bF_buf4), .Y(_8968_) );
	OAI21X1 OAI21X1_3790 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_8847__bF_buf7), .C(_8968_), .Y(_8969_) );
	AOI21X1 AOI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_8967_), .C(_7303__bF_buf4_bF_buf3), .Y(_8970_) );
	OAI21X1 OAI21X1_3791 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_7842_), .C(_8970_), .Y(_8971_) );
	AOI21X1 AOI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .B(_8969_), .C(rst_bF_buf18), .Y(_6709__22_) );
	INVX1 INVX1_1561 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_23_), .Y(_8972_) );
	AOI21X1 AOI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf6), .B(_8972_), .C(_7304__bF_buf3), .Y(_8973_) );
	OAI21X1 OAI21X1_3792 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf3), .B(_8847__bF_buf5), .C(_8973_), .Y(_8974_) );
	AOI21X1 AOI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_8972_), .C(_7303__bF_buf3_bF_buf3), .Y(_8975_) );
	OAI21X1 OAI21X1_3793 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_7857_), .C(_8975_), .Y(_8976_) );
	AOI21X1 AOI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_8976_), .B(_8974_), .C(rst_bF_buf17), .Y(_6709__23_) );
	INVX1 INVX1_1562 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_24_), .Y(_8977_) );
	AOI21X1 AOI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf4), .B(_8977_), .C(_7304__bF_buf2), .Y(_8978_) );
	OAI21X1 OAI21X1_3794 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_8847__bF_buf3), .C(_8978_), .Y(_8979_) );
	AOI21X1 AOI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_8977_), .C(_7303__bF_buf2), .Y(_8980_) );
	OAI21X1 OAI21X1_3795 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_7865_), .C(_8980_), .Y(_8981_) );
	AOI21X1 AOI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_8981_), .B(_8979_), .C(rst_bF_buf16), .Y(_6709__24_) );
	INVX1 INVX1_1563 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_25_), .Y(_8982_) );
	AOI21X1 AOI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf2), .B(_8982_), .C(_7304__bF_buf1), .Y(_8983_) );
	OAI21X1 OAI21X1_3796 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf1), .B(_8847__bF_buf1), .C(_8983_), .Y(_8984_) );
	AOI21X1 AOI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_8982_), .C(_7303__bF_buf1), .Y(_8985_) );
	OAI21X1 OAI21X1_3797 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_7881_), .C(_8985_), .Y(_8986_) );
	AOI21X1 AOI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_8986_), .B(_8984_), .C(rst_bF_buf15), .Y(_6709__25_) );
	OAI21X1 OAI21X1_3798 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_7424__bF_buf2), .C(csr_gpr_iu_csr_mepc_26_), .Y(_8987_) );
	OAI21X1 OAI21X1_3799 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_7890_), .C(_8987_), .Y(_8988_) );
	OAI21X1 OAI21X1_3800 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf1), .C(_8988_), .Y(_8989_) );
	AOI21X1 AOI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_8846__bF_buf2), .B(_7405_), .C(_7304__bF_buf0), .Y(_8990_) );
	OAI21X1 OAI21X1_3801 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_26_), .B(_8846__bF_buf1), .C(_8990_), .Y(_8991_) );
	AOI21X1 AOI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_8989_), .B(_8991_), .C(rst_bF_buf14), .Y(_6709__26_) );
	NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_8616__bF_buf7), .B(_7897_), .Y(_8992_) );
	OAI21X1 OAI21X1_3802 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_27_), .B(_8616__bF_buf6), .C(_8992_), .Y(_8993_) );
	NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_7555_), .B(_8847__bF_buf0), .Y(_8994_) );
	INVX1 INVX1_1564 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_27_), .Y(_8995_) );
	OAI21X1 OAI21X1_3803 ( .gnd(gnd), .vdd(vdd), .A(_8995_), .B(_8893_), .C(_7303__bF_buf0), .Y(_8996_) );
	OAI21X1 OAI21X1_3804 ( .gnd(gnd), .vdd(vdd), .A(_8996_), .B(_8994_), .C(_6879__bF_buf16), .Y(_8997_) );
	AOI21X1 AOI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_8993_), .B(_7304__bF_buf14_bF_buf3), .C(_8997_), .Y(_6709__27_) );
	NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_8616__bF_buf5), .B(_7907_), .Y(_8998_) );
	OAI21X1 OAI21X1_3805 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_28_), .B(_8616__bF_buf4), .C(_8998_), .Y(_8999_) );
	NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_8847__bF_buf7), .Y(_9000_) );
	INVX1 INVX1_1565 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_28_), .Y(_9001_) );
	OAI21X1 OAI21X1_3806 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8893_), .C(_7303__bF_buf14_bF_buf2), .Y(_9002_) );
	OAI21X1 OAI21X1_3807 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_9000_), .C(_6879__bF_buf15), .Y(_9003_) );
	AOI21X1 AOI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_8999_), .B(_7304__bF_buf13_bF_buf3), .C(_9003_), .Y(_6709__28_) );
	INVX1 INVX1_1566 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_29_), .Y(_9004_) );
	AOI21X1 AOI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf6), .B(_9004_), .C(_7304__bF_buf12_bF_buf3), .Y(_9005_) );
	OAI21X1 OAI21X1_3808 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf1), .B(_8847__bF_buf5), .C(_9005_), .Y(_9006_) );
	AOI21X1 AOI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_9004_), .C(_7303__bF_buf13_bF_buf2), .Y(_9007_) );
	OAI21X1 OAI21X1_3809 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf6), .B(_7928_), .C(_9007_), .Y(_9008_) );
	AOI21X1 AOI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_9008_), .B(_9006_), .C(rst_bF_buf13), .Y(_6709__29_) );
	INVX1 INVX1_1567 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_30_), .Y(_9009_) );
	AOI21X1 AOI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf4), .B(_9009_), .C(_7304__bF_buf11_bF_buf3), .Y(_9010_) );
	OAI21X1 OAI21X1_3810 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_8847__bF_buf3), .C(_9010_), .Y(_9011_) );
	AOI21X1 AOI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf5), .B(_9009_), .C(_7303__bF_buf12_bF_buf2), .Y(_9012_) );
	OAI21X1 OAI21X1_3811 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf4), .B(_7941_), .C(_9012_), .Y(_9013_) );
	AOI21X1 AOI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_9013_), .B(_9011_), .C(rst_bF_buf12), .Y(_6709__30_) );
	INVX1 INVX1_1568 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_31_), .Y(_9014_) );
	AOI21X1 AOI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf2), .B(_9014_), .C(_7304__bF_buf10_bF_buf3), .Y(_9015_) );
	OAI21X1 OAI21X1_3812 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf3), .B(_8847__bF_buf1), .C(_9015_), .Y(_9016_) );
	AOI21X1 AOI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf3), .B(_9014_), .C(_7303__bF_buf11_bF_buf2), .Y(_9017_) );
	OAI21X1 OAI21X1_3813 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf2), .B(_7949_), .C(_9017_), .Y(_9018_) );
	AOI21X1 AOI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_9018_), .B(_9016_), .C(rst_bF_buf11), .Y(_6709__31_) );
	NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .B(_8060_), .Y(_9019_) );
	NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf5), .B(_7304__bF_buf9_bF_buf3), .Y(_9020_) );
	INVX8 INVX8_80 ( .gnd(gnd), .vdd(vdd), .A(_9020__bF_buf3), .Y(_9021_) );
	OAI21X1 OAI21X1_3814 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf4), .B(_7304__bF_buf8_bF_buf3), .C(csr_gpr_iu_csr_mtvec_0_), .Y(_9022_) );
	OAI21X1 OAI21X1_3815 ( .gnd(gnd), .vdd(vdd), .A(_7324_), .B(_9021__bF_buf4), .C(_9022_), .Y(_9023_) );
	AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_6879__bF_buf14), .Y(_6723__0_) );
	OAI21X1 OAI21X1_3816 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf3), .B(_7304__bF_buf7_bF_buf3), .C(csr_gpr_iu_csr_mtvec_1_), .Y(_9024_) );
	OAI21X1 OAI21X1_3817 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_9021__bF_buf3), .C(_9024_), .Y(_9025_) );
	AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_9025_), .B(_6879__bF_buf13), .Y(_6723__1_) );
	OAI21X1 OAI21X1_3818 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf2), .B(_7304__bF_buf6_bF_buf3), .C(csr_gpr_iu_csr_mtvec_2_), .Y(_9026_) );
	NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_9020__bF_buf2), .Y(_9027_) );
	AOI21X1 AOI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(_9026_), .C(rst_bF_buf10), .Y(_6723__2_) );
	INVX1 INVX1_1569 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_3_), .Y(_9028_) );
	OAI21X1 OAI21X1_3819 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf1), .B(_7304__bF_buf5), .C(_9028_), .Y(_9029_) );
	OAI21X1 OAI21X1_3820 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_9021__bF_buf2), .C(_9029_), .Y(_9030_) );
	NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf9), .B(_9030_), .Y(_6723__3_) );
	OAI21X1 OAI21X1_3821 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf0), .B(_7304__bF_buf4), .C(csr_gpr_iu_csr_mtvec_4_), .Y(_9031_) );
	NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_9020__bF_buf1), .Y(_9032_) );
	AOI21X1 AOI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_9032_), .B(_9031_), .C(rst_bF_buf8), .Y(_6723__4_) );
	OAI21X1 OAI21X1_3822 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf5), .B(_7304__bF_buf3), .C(csr_gpr_iu_csr_mtvec_5_), .Y(_9033_) );
	NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_9020__bF_buf0), .Y(_9034_) );
	AOI21X1 AOI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9033_), .C(rst_bF_buf7), .Y(_6723__5_) );
	OAI21X1 OAI21X1_3823 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf4), .B(_7304__bF_buf2), .C(csr_gpr_iu_csr_mtvec_6_), .Y(_9035_) );
	NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_9020__bF_buf3), .Y(_9036_) );
	AOI21X1 AOI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_9036_), .B(_9035_), .C(rst_bF_buf6), .Y(_6723__6_) );
	OAI21X1 OAI21X1_3824 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf3), .B(_7304__bF_buf1), .C(csr_gpr_iu_csr_mtvec_7_), .Y(_9037_) );
	NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_9020__bF_buf2), .Y(_9038_) );
	AOI21X1 AOI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_9038_), .B(_9037_), .C(rst_bF_buf5), .Y(_6723__7_) );
	OAI21X1 OAI21X1_3825 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf2), .B(_7304__bF_buf0), .C(csr_gpr_iu_csr_mtvec_8_), .Y(_9039_) );
	NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_9020__bF_buf1), .Y(_9040_) );
	AOI21X1 AOI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_9039_), .C(rst_bF_buf4), .Y(_6723__8_) );
	OAI21X1 OAI21X1_3826 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf1), .B(_7304__bF_buf14_bF_buf2), .C(csr_gpr_iu_csr_mtvec_9_), .Y(_9041_) );
	NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_9020__bF_buf0), .Y(_9042_) );
	AOI21X1 AOI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_9041_), .C(rst_bF_buf3), .Y(_6723__9_) );
	OAI21X1 OAI21X1_3827 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf0), .B(_7304__bF_buf13_bF_buf2), .C(csr_gpr_iu_csr_mtvec_10_), .Y(_9043_) );
	NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_9020__bF_buf3), .Y(_9044_) );
	AOI21X1 AOI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .B(_9043_), .C(rst_bF_buf2), .Y(_6723__10_) );
	OAI21X1 OAI21X1_3828 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf5), .B(_7304__bF_buf12_bF_buf2), .C(csr_gpr_iu_csr_mtvec_11_), .Y(_9045_) );
	NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .B(_9020__bF_buf2), .Y(_9046_) );
	AOI21X1 AOI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_9046_), .B(_9045_), .C(rst_bF_buf1), .Y(_6723__11_) );
	OAI21X1 OAI21X1_3829 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf4), .B(_7304__bF_buf11_bF_buf2), .C(csr_gpr_iu_csr_mtvec_12_), .Y(_9047_) );
	NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_9020__bF_buf1), .Y(_9048_) );
	AOI21X1 AOI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_9048_), .B(_9047_), .C(rst_bF_buf0), .Y(_6723__12_) );
	INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_13_), .Y(_9049_) );
	OAI21X1 OAI21X1_3830 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf1), .B(_9021__bF_buf1), .C(_6879__bF_buf12), .Y(_9050_) );
	AOI21X1 AOI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_9049_), .B(_9021__bF_buf0), .C(_9050_), .Y(_6723__13_) );
	OAI21X1 OAI21X1_3831 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf3), .B(_7304__bF_buf10_bF_buf2), .C(csr_gpr_iu_csr_mtvec_14_), .Y(_9051_) );
	NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_9020__bF_buf0), .Y(_9052_) );
	AOI21X1 AOI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_9052_), .B(_9051_), .C(rst_bF_buf70), .Y(_6723__14_) );
	INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_15_), .Y(_9053_) );
	OAI21X1 OAI21X1_3832 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf2), .B(_9021__bF_buf4), .C(_6879__bF_buf11), .Y(_9054_) );
	AOI21X1 AOI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_9021__bF_buf3), .C(_9054_), .Y(_6723__15_) );
	OAI21X1 OAI21X1_3833 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf2), .B(_7304__bF_buf9_bF_buf2), .C(csr_gpr_iu_csr_mtvec_16_), .Y(_9055_) );
	NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_9020__bF_buf3), .Y(_9056_) );
	AOI21X1 AOI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_9056_), .B(_9055_), .C(rst_bF_buf69), .Y(_6723__16_) );
	INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_17_), .Y(_9057_) );
	OAI21X1 OAI21X1_3834 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf3), .B(_9021__bF_buf2), .C(_6879__bF_buf10), .Y(_9058_) );
	AOI21X1 AOI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_9021__bF_buf1), .C(_9058_), .Y(_6723__17_) );
	OAI21X1 OAI21X1_3835 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf1), .B(_7304__bF_buf8_bF_buf2), .C(csr_gpr_iu_csr_mtvec_18_), .Y(_9059_) );
	OAI21X1 OAI21X1_3836 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_9021__bF_buf0), .C(_9059_), .Y(_9060_) );
	AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_9060_), .B(_6879__bF_buf9), .Y(_6723__18_) );
	INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_19_), .Y(_9061_) );
	OAI21X1 OAI21X1_3837 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf0), .B(_9021__bF_buf4), .C(_6879__bF_buf8), .Y(_9062_) );
	AOI21X1 AOI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_9021__bF_buf3), .C(_9062_), .Y(_6723__19_) );
	OAI21X1 OAI21X1_3838 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf0), .B(_7304__bF_buf7_bF_buf2), .C(csr_gpr_iu_csr_mtvec_20_), .Y(_9063_) );
	OAI21X1 OAI21X1_3839 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_9021__bF_buf2), .C(_9063_), .Y(_9064_) );
	AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_9064_), .B(_6879__bF_buf7), .Y(_6723__20_) );
	INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_21_), .Y(_9065_) );
	OAI21X1 OAI21X1_3840 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf0), .B(_9021__bF_buf1), .C(_6879__bF_buf6), .Y(_9066_) );
	AOI21X1 AOI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9021__bF_buf0), .C(_9066_), .Y(_6723__21_) );
	NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_9020__bF_buf2), .Y(_9067_) );
	OAI21X1 OAI21X1_3841 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_22_), .B(_9020__bF_buf1), .C(_9067_), .Y(_9068_) );
	NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf68), .B(_9068_), .Y(_6723__22_) );
	INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_23_), .Y(_9069_) );
	OAI21X1 OAI21X1_3842 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf2), .B(_9021__bF_buf4), .C(_6879__bF_buf5), .Y(_9070_) );
	AOI21X1 AOI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_9069_), .B(_9021__bF_buf3), .C(_9070_), .Y(_6723__23_) );
	OAI21X1 OAI21X1_3843 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf5), .B(_7304__bF_buf6_bF_buf2), .C(csr_gpr_iu_csr_mtvec_24_), .Y(_9071_) );
	NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_9020__bF_buf0), .Y(_9072_) );
	AOI21X1 AOI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(_9071_), .C(rst_bF_buf67), .Y(_6723__24_) );
	INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_25_), .Y(_9073_) );
	OAI21X1 OAI21X1_3844 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf0), .B(_9021__bF_buf2), .C(_6879__bF_buf4), .Y(_9074_) );
	AOI21X1 AOI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_9073_), .B(_9021__bF_buf1), .C(_9074_), .Y(_6723__25_) );
	OAI21X1 OAI21X1_3845 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf4), .B(_7304__bF_buf5), .C(csr_gpr_iu_csr_mtvec_26_), .Y(_9075_) );
	OAI21X1 OAI21X1_3846 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_9021__bF_buf0), .C(_9075_), .Y(_9076_) );
	AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(_6879__bF_buf3), .Y(_6723__26_) );
	INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_27_), .Y(_9077_) );
	OAI21X1 OAI21X1_3847 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf1), .B(_9021__bF_buf4), .C(_6879__bF_buf2), .Y(_9078_) );
	AOI21X1 AOI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_9077_), .B(_9021__bF_buf3), .C(_9078_), .Y(_6723__27_) );
	OAI21X1 OAI21X1_3848 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf3), .B(_7304__bF_buf4), .C(csr_gpr_iu_csr_mtvec_28_), .Y(_9079_) );
	NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_9020__bF_buf3), .Y(_9080_) );
	AOI21X1 AOI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_9080_), .B(_9079_), .C(rst_bF_buf66), .Y(_6723__28_) );
	INVX1 INVX1_1570 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_29_), .Y(_9081_) );
	OAI21X1 OAI21X1_3849 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf0), .B(_9021__bF_buf2), .C(_6879__bF_buf1), .Y(_9082_) );
	AOI21X1 AOI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_9081_), .B(_9021__bF_buf1), .C(_9082_), .Y(_6723__29_) );
	OAI21X1 OAI21X1_3850 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf2), .B(_7304__bF_buf3), .C(csr_gpr_iu_csr_mtvec_30_), .Y(_9083_) );
	NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_9020__bF_buf2), .Y(_9084_) );
	AOI21X1 AOI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_9083_), .C(rst_bF_buf65), .Y(_6723__30_) );
	INVX1 INVX1_1571 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_31_), .Y(_9085_) );
	OAI21X1 OAI21X1_3851 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf2), .B(_9021__bF_buf0), .C(_6879__bF_buf0), .Y(_9086_) );
	AOI21X1 AOI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_9085_), .B(_9021__bF_buf4), .C(_9086_), .Y(_6723__31_) );
	NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_8057_), .Y(_9087_) );
	OAI21X1 OAI21X1_3852 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .B(_7308_), .C(_9087_), .Y(_9088_) );
	INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .Y(_9089_) );
	OAI21X1 OAI21X1_3853 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_9089_), .C(csr_gpr_iu_csr_sie), .Y(_9090_) );
	OAI21X1 OAI21X1_3854 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_9088_), .C(_9090_), .Y(_9091_) );
	NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf2), .B(_9091_), .Y(_9092_) );
	INVX1 INVX1_1572 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_ret), .Y(_9093_) );
	NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_9093_), .B(_6930__bF_buf0), .Y(_9094_) );
	INVX8 INVX8_81 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf5), .Y(_9095_) );
	NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sie), .B(_7594__bF_buf6), .C(_9095__bF_buf4), .Y(_9096_) );
	INVX4 INVX4_20 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf3), .Y(_9097_) );
	NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .B(_9097_), .Y(_9098_) );
	MUX2X1 MUX2X1_159 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spie), .B(csr_gpr_iu_csr_sie), .S(_9098__bF_buf4), .Y(_9099_) );
	OAI21X1 OAI21X1_3855 ( .gnd(gnd), .vdd(vdd), .A(_9095__bF_buf3), .B(_9099_), .C(_9096_), .Y(_9100_) );
	OAI21X1 OAI21X1_3856 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf5), .C(_9100_), .Y(_9101_) );
	AOI21X1 AOI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_9101_), .B(_9092_), .C(rst_bF_buf64), .Y(_6743_) );
	INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mie), .Y(_9102_) );
	INVX1 INVX1_1573 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .Y(_9103_) );
	NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_9103_), .Y(_9104_) );
	INVX8 INVX8_82 ( .gnd(gnd), .vdd(vdd), .A(_9104_), .Y(_9105_) );
	OAI21X1 OAI21X1_3857 ( .gnd(gnd), .vdd(vdd), .A(_9105__bF_buf4), .B(_9095__bF_buf2), .C(_9102_), .Y(_9106_) );
	INVX1 INVX1_1574 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpie), .Y(_9107_) );
	NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_9104_), .C(_9094__bF_buf4), .Y(_9108_) );
	NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf1), .B(_9108_), .C(_9106_), .Y(_9109_) );
	NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_8111__bF_buf3), .Y(_9110_) );
	NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_9110__bF_buf3), .Y(_9111_) );
	OAI21X1 OAI21X1_3858 ( .gnd(gnd), .vdd(vdd), .A(_9102_), .B(_9110__bF_buf2), .C(_9111_), .Y(_9112_) );
	OAI21X1 OAI21X1_3859 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf2), .B(_9112_), .C(_6879__bF_buf42), .Y(_9113_) );
	AOI21X1 AOI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_7304__bF_buf1), .B(_9109_), .C(_9113_), .Y(_6711_) );
	NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_9110__bF_buf1), .Y(_9114_) );
	OAI21X1 OAI21X1_3860 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spie), .B(_9110__bF_buf0), .C(_9114_), .Y(_9115_) );
	NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spie), .B(_7428__bF_buf2), .Y(_9116_) );
	AOI21X1 AOI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_9102_), .B(_7428__bF_buf1), .C(_9116_), .Y(_9117_) );
	OAI21X1 OAI21X1_3861 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9_bF_buf2), .B(_9117_), .C(_6879__bF_buf41), .Y(_9118_) );
	AOI21X1 AOI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_9115_), .B(_7303__bF_buf8_bF_buf2), .C(_9118_), .Y(_6744_) );
	NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_9110__bF_buf3), .Y(_9119_) );
	OAI21X1 OAI21X1_3862 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpie), .B(_9110__bF_buf2), .C(_9119_), .Y(_9120_) );
	MUX2X1 MUX2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_9102_), .B(_9107_), .S(_8616__bF_buf3), .Y(_9121_) );
	OAI21X1 OAI21X1_3863 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf7_bF_buf2), .B(_9121_), .C(_6879__bF_buf40), .Y(_9122_) );
	AOI21X1 AOI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(_7303__bF_buf6_bF_buf2), .C(_9122_), .Y(_6713_) );
	INVX1 INVX1_1575 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spp), .Y(_9123_) );
	OAI21X1 OAI21X1_3864 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_9089_), .C(_9123_), .Y(_9124_) );
	OAI21X1 OAI21X1_3865 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_9088_), .C(_9124_), .Y(_9125_) );
	NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf2), .B(biu_mmu_msu_1_), .Y(_9126_) );
	MUX2X1 MUX2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9123_), .S(_7428__bF_buf0), .Y(_9127_) );
	OAI21X1 OAI21X1_3866 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf5_bF_buf2), .B(_9127_), .C(_6879__bF_buf39), .Y(_9128_) );
	AOI21X1 AOI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_9125_), .B(_7303__bF_buf4_bF_buf2), .C(_9128_), .Y(_6745_) );
	NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_9110__bF_buf1), .Y(_9129_) );
	OAI21X1 OAI21X1_3867 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_0_), .B(_9110__bF_buf0), .C(_9129_), .Y(_9130_) );
	INVX1 INVX1_1576 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_0_), .Y(_9131_) );
	MUX2X1 MUX2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_9131_), .S(_8616__bF_buf2), .Y(_9132_) );
	OAI21X1 OAI21X1_3868 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf3_bF_buf2), .B(_9132_), .C(_6879__bF_buf38), .Y(_9133_) );
	AOI21X1 AOI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_9130_), .B(_7303__bF_buf2), .C(_9133_), .Y(_6714__0_) );
	NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_9110__bF_buf3), .Y(_9134_) );
	OAI21X1 OAI21X1_3869 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_1_), .B(_9110__bF_buf2), .C(_9134_), .Y(_9135_) );
	NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_1_), .B(_8616__bF_buf1), .Y(_9136_) );
	AOI21X1 AOI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_9103_), .B(_8616__bF_buf0), .C(_9136_), .Y(_9137_) );
	OAI21X1 OAI21X1_3870 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf1), .B(_9137_), .C(_6879__bF_buf37), .Y(_9138_) );
	AOI21X1 AOI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_9135_), .B(_7303__bF_buf0), .C(_9138_), .Y(_6714__1_) );
	INVX1 INVX1_1577 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mprv), .Y(_9139_) );
	NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf14_bF_buf1), .B(_9110__bF_buf1), .Y(_9140_) );
	OAI21X1 OAI21X1_3871 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf2), .B(_9140_), .C(_6879__bF_buf36), .Y(_9141_) );
	AOI21X1 AOI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(_9140_), .C(_9141_), .Y(_6715_) );
	MUX2X1 MUX2X1_163 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_tvm), .B(addr_csr_20_), .S(_9140_), .Y(_9142_) );
	NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf63), .B(_9142_), .Y(_6755_) );
	MUX2X1 MUX2X1_164 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_tsr), .B(addr_csr_22_), .S(_9140_), .Y(_9143_) );
	NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf62), .B(_9143_), .Y(_6754_) );
	NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_7309__bF_buf1), .Y(_9144_) );
	OAI21X1 OAI21X1_3872 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf0), .B(_9144_), .C(_7303__bF_buf13_bF_buf1), .Y(_9145_) );
	MUX2X1 MUX2X1_165 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_sum), .B(addr_csr_18_), .S(_9145_), .Y(_9146_) );
	NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf61), .B(_9146_), .Y(_6753_) );
	INVX1 INVX1_1578 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_mxr), .Y(_9147_) );
	OAI21X1 OAI21X1_3873 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf3), .B(_9145_), .C(_6879__bF_buf35), .Y(_9148_) );
	AOI21X1 AOI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_9145_), .C(_9148_), .Y(_6724_) );
	NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7424__bF_buf1), .Y(_9149_) );
	OAI21X1 OAI21X1_3874 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf12_bF_buf1), .B(_9095__bF_buf1), .C(_9097_), .Y(_9150_) );
	NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_9149__bF_buf4), .B(_9150_), .Y(_9151_) );
	OAI21X1 OAI21X1_3875 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_6930__bF_buf4), .C(_9094__bF_buf3), .Y(_9152_) );
	NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spp), .B(_9098__bF_buf3), .Y(_9153_) );
	OAI21X1 OAI21X1_3876 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .B(_9105__bF_buf3), .C(_9153_), .Y(_9154_) );
	NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_9152_), .Y(_9155_) );
	OAI21X1 OAI21X1_3877 ( .gnd(gnd), .vdd(vdd), .A(_9155_), .B(_9151_), .C(_6879__bF_buf34), .Y(_6719__0_) );
	OAI21X1 OAI21X1_3878 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(csr_gpr_iu_csr_mpp_1_), .C(_9094__bF_buf2), .Y(_9156_) );
	OAI21X1 OAI21X1_3879 ( .gnd(gnd), .vdd(vdd), .A(_7428__bF_buf8), .B(_9094__bF_buf1), .C(_9156_), .Y(_9157_) );
	OAI22X1 OAI22X1_745 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .B(_9149__bF_buf3), .C(_7303__bF_buf11_bF_buf1), .D(_9157_), .Y(_9158_) );
	NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_6879__bF_buf33), .B(_9158_), .Y(_6719__1_) );
	NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_8113_), .Y(_9159_) );
	NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_9159_), .Y(_9160_) );
	NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_9160_), .B(_7308_), .Y(_9161_) );
	NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf4), .B(_7304__bF_buf0), .Y(_9162_) );
	NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_7324_), .B(_9162__bF_buf3), .Y(_9163_) );
	OAI21X1 OAI21X1_3880 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_12_), .B(_9162__bF_buf2), .C(_9163_), .Y(_9164_) );
	NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf60), .B(_9164_), .Y(_6738__0_) );
	NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_9162__bF_buf1), .Y(_9165_) );
	OAI21X1 OAI21X1_3881 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_13_), .B(_9162__bF_buf0), .C(_9165_), .Y(_9166_) );
	NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf59), .B(_9166_), .Y(_6738__1_) );
	OAI21X1 OAI21X1_3882 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf3), .B(_7304__bF_buf14_bF_buf1), .C(biu_mmu_ag0_14_), .Y(_9167_) );
	NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_9162__bF_buf3), .Y(_9168_) );
	AOI21X1 AOI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_9168_), .B(_9167_), .C(rst_bF_buf58), .Y(_6738__2_) );
	NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_6895_), .B(_9162__bF_buf2), .Y(_9169_) );
	OAI21X1 OAI21X1_3883 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_15_), .B(_9162__bF_buf1), .C(_9169_), .Y(_9170_) );
	NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf57), .B(_9170_), .Y(_6738__3_) );
	OAI21X1 OAI21X1_3884 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf2), .B(_7304__bF_buf13_bF_buf1), .C(biu_mmu_ag0_16_), .Y(_9171_) );
	NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_9162__bF_buf0), .Y(_9172_) );
	AOI21X1 AOI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_9172_), .B(_9171_), .C(rst_bF_buf56), .Y(_6738__4_) );
	NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_9162__bF_buf3), .Y(_9173_) );
	OAI21X1 OAI21X1_3885 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_17_), .B(_9162__bF_buf2), .C(_9173_), .Y(_9174_) );
	NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf55), .B(_9174_), .Y(_6738__5_) );
	INVX8 INVX8_83 ( .gnd(gnd), .vdd(vdd), .A(_9162__bF_buf1), .Y(_9175_) );
	OAI21X1 OAI21X1_3886 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf1), .B(_7304__bF_buf12_bF_buf1), .C(biu_mmu_ag0_18_), .Y(_9176_) );
	OAI21X1 OAI21X1_3887 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_9175__bF_buf4), .C(_9176_), .Y(_9177_) );
	AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_6879__bF_buf32), .Y(_6738__6_) );
	NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_9162__bF_buf0), .Y(_9178_) );
	OAI21X1 OAI21X1_3888 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_19_), .B(_9162__bF_buf3), .C(_9178_), .Y(_9179_) );
	NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf54), .B(_9179_), .Y(_6738__7_) );
	OAI21X1 OAI21X1_3889 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf0), .B(_7304__bF_buf11_bF_buf1), .C(biu_mmu_ag0_20_), .Y(_9180_) );
	OAI21X1 OAI21X1_3890 ( .gnd(gnd), .vdd(vdd), .A(_6927_), .B(_9175__bF_buf3), .C(_9180_), .Y(_9181_) );
	AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_9181_), .B(_6879__bF_buf31), .Y(_6738__8_) );
	NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_9162__bF_buf2), .Y(_9182_) );
	OAI21X1 OAI21X1_3891 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_21_), .B(_9162__bF_buf1), .C(_9182_), .Y(_9183_) );
	NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf53), .B(_9183_), .Y(_6738__9_) );
	NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_9162__bF_buf0), .Y(_9184_) );
	OAI21X1 OAI21X1_3892 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_22_), .B(_9162__bF_buf3), .C(_9184_), .Y(_9185_) );
	NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf52), .B(_9185_), .Y(_6738__10_) );
	NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_9162__bF_buf2), .Y(_9186_) );
	OAI21X1 OAI21X1_3893 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_23_), .B(_9162__bF_buf1), .C(_9186_), .Y(_9187_) );
	NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf51), .B(_9187_), .Y(_6738__11_) );
	INVX1 INVX1_1579 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_24_), .Y(_9188_) );
	OAI21X1 OAI21X1_3894 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf4), .B(_7304__bF_buf10_bF_buf1), .C(_9188_), .Y(_9189_) );
	OAI21X1 OAI21X1_3895 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_9175__bF_buf2), .C(_9189_), .Y(_9190_) );
	NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf50), .B(_9190_), .Y(_6738__12_) );
	INVX1 INVX1_1580 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_25_), .Y(_9191_) );
	OAI21X1 OAI21X1_3896 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf0), .B(_9175__bF_buf1), .C(_6879__bF_buf30), .Y(_9192_) );
	AOI21X1 AOI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_9175__bF_buf0), .C(_9192_), .Y(_6738__13_) );
	OAI21X1 OAI21X1_3897 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf3), .B(_7304__bF_buf9_bF_buf1), .C(biu_mmu_ag0_26_), .Y(_9193_) );
	NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_9162__bF_buf0), .Y(_9194_) );
	AOI21X1 AOI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_9193_), .C(rst_bF_buf49), .Y(_6738__14_) );
	INVX1 INVX1_1581 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_27_), .Y(_9195_) );
	OAI21X1 OAI21X1_3898 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf1), .B(_9175__bF_buf4), .C(_6879__bF_buf29), .Y(_9196_) );
	AOI21X1 AOI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_9195_), .B(_9175__bF_buf3), .C(_9196_), .Y(_6738__15_) );
	OAI21X1 OAI21X1_3899 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf2), .B(_7304__bF_buf8_bF_buf1), .C(biu_mmu_ag0_28_), .Y(_9197_) );
	OAI21X1 OAI21X1_3900 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_9175__bF_buf2), .C(_9197_), .Y(_9198_) );
	AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(_6879__bF_buf28), .Y(_6738__16_) );
	INVX1 INVX1_1582 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_29_), .Y(_9199_) );
	OAI21X1 OAI21X1_3901 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf1), .B(_9175__bF_buf1), .C(_6879__bF_buf27), .Y(_9200_) );
	AOI21X1 AOI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_9199_), .B(_9175__bF_buf0), .C(_9200_), .Y(_6738__17_) );
	OAI21X1 OAI21X1_3902 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf1), .B(_7304__bF_buf7_bF_buf1), .C(biu_mmu_ag0_30_), .Y(_9201_) );
	OAI21X1 OAI21X1_3903 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_9175__bF_buf4), .C(_9201_), .Y(_9202_) );
	AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(_6879__bF_buf26), .Y(_6738__18_) );
	INVX1 INVX1_1583 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_31_), .Y(_9203_) );
	OAI21X1 OAI21X1_3904 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf2), .B(_9175__bF_buf3), .C(_6879__bF_buf25), .Y(_9204_) );
	AOI21X1 AOI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_9175__bF_buf2), .C(_9204_), .Y(_6738__19_) );
	INVX1 INVX1_1584 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_32_), .Y(_9205_) );
	OAI21X1 OAI21X1_3905 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf0), .B(_7304__bF_buf6_bF_buf1), .C(_9205_), .Y(_9206_) );
	OAI21X1 OAI21X1_3906 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_9175__bF_buf1), .C(_9206_), .Y(_9207_) );
	NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf48), .B(_9207_), .Y(_6738__20_) );
	INVX1 INVX1_1585 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_33_), .Y(_9208_) );
	OAI21X1 OAI21X1_3907 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf3), .B(_9175__bF_buf0), .C(_6879__bF_buf24), .Y(_9209_) );
	AOI21X1 AOI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_9175__bF_buf4), .C(_9209_), .Y(_6738__21_) );
	INVX1 INVX1_1586 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_22_), .Y(_9210_) );
	OAI21X1 OAI21X1_3908 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf4), .B(_7304__bF_buf5), .C(_9210_), .Y(_9211_) );
	OAI21X1 OAI21X1_3909 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_9175__bF_buf3), .C(_9211_), .Y(_9212_) );
	NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf47), .B(_9212_), .Y(_6738__22_) );
	INVX1 INVX1_1587 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_23_), .Y(_9213_) );
	OAI21X1 OAI21X1_3910 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf1), .B(_9175__bF_buf2), .C(_6879__bF_buf23), .Y(_9214_) );
	AOI21X1 AOI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_9175__bF_buf1), .C(_9214_), .Y(_6738__23_) );
	OAI21X1 OAI21X1_3911 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf3), .B(_7304__bF_buf4), .C(biu_mmu_satp_24_), .Y(_9215_) );
	OAI21X1 OAI21X1_3912 ( .gnd(gnd), .vdd(vdd), .A(_7399_), .B(_9175__bF_buf0), .C(_9215_), .Y(_9216_) );
	AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(_6879__bF_buf22), .Y(_6738__24_) );
	INVX1 INVX1_1588 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_25_), .Y(_9217_) );
	OAI21X1 OAI21X1_3913 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf3), .B(_9175__bF_buf4), .C(_6879__bF_buf21), .Y(_9218_) );
	AOI21X1 AOI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_9175__bF_buf3), .C(_9218_), .Y(_6738__25_) );
	NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_9162__bF_buf3), .Y(_9219_) );
	OAI21X1 OAI21X1_3914 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_26_), .B(_9162__bF_buf2), .C(_9219_), .Y(_9220_) );
	NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf46), .B(_9220_), .Y(_6738__26_) );
	INVX1 INVX1_1589 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_27_), .Y(_9221_) );
	OAI21X1 OAI21X1_3915 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf0), .B(_9175__bF_buf2), .C(_6879__bF_buf20), .Y(_9222_) );
	AOI21X1 AOI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_9221_), .B(_9175__bF_buf1), .C(_9222_), .Y(_6738__27_) );
	OAI21X1 OAI21X1_3916 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf2), .B(_7304__bF_buf3), .C(biu_mmu_satp_28_), .Y(_9223_) );
	OAI21X1 OAI21X1_3917 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_9175__bF_buf0), .C(_9223_), .Y(_9224_) );
	AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_9224_), .B(_6879__bF_buf19), .Y(_6738__28_) );
	INVX1 INVX1_1590 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_29_), .Y(_9225_) );
	OAI21X1 OAI21X1_3918 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf3), .B(_9175__bF_buf4), .C(_6879__bF_buf18), .Y(_9226_) );
	AOI21X1 AOI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_9225_), .B(_9175__bF_buf3), .C(_9226_), .Y(_6738__29_) );
	OAI21X1 OAI21X1_3919 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf1), .B(_7304__bF_buf2), .C(biu_mmu_satp_30_), .Y(_9227_) );
	NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_9162__bF_buf1), .Y(_9228_) );
	AOI21X1 AOI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_9228_), .B(_9227_), .C(rst_bF_buf45), .Y(_6738__30_) );
	INVX1 INVX1_1591 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_31_), .Y(_9229_) );
	OAI21X1 OAI21X1_3920 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf1), .B(_9175__bF_buf2), .C(_6879__bF_buf17), .Y(_9230_) );
	AOI21X1 AOI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_9175__bF_buf1), .C(_9230_), .Y(_6738__31_) );
	OAI21X1 OAI21X1_3921 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_7582_), .C(_7957_), .Y(_9231_) );
	NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .B(_9231_), .C(_8116_), .Y(_9232_) );
	INVX1 INVX1_1592 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf2), .Y(_9233_) );
	INVX8 INVX8_84 ( .gnd(gnd), .vdd(vdd), .A(_9161__bF_buf0), .Y(_9234_) );
	OAI21X1 OAI21X1_3922 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_9089_), .C(_9019__bF_buf1), .Y(_9235_) );
	NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .B(_9234__bF_buf3), .Y(_9236_) );
	NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_8062__bF_buf0), .Y(_9237_) );
	NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_9233_), .B(_9236_), .C(_9237_), .Y(_9238_) );
	OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_9238_), .B(_9232_), .Y(_9239_) );
	OAI21X1 OAI21X1_3923 ( .gnd(gnd), .vdd(vdd), .A(_8161_), .B(_8112_), .C(_7317_), .Y(_9240_) );
	OAI21X1 OAI21X1_3924 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_8325_), .C(_8278_), .Y(_9241_) );
	NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_8486__bF_buf1), .B(_9241_), .C(_8554_), .Y(_9242_) );
	OAI21X1 OAI21X1_3925 ( .gnd(gnd), .vdd(vdd), .A(_8231_), .B(_8161_), .C(_8115_), .Y(_9243_) );
	NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .B(_8326_), .C(_9243_), .Y(_9244_) );
	NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_9242_), .B(_9244_), .Y(_9245_) );
	NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_8847__bF_buf0), .B(_9240_), .C(_9245_), .Y(_9246_) );
	NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9246_), .Y(_9247_) );
	NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_9247_), .Y(_9248_) );
	OAI21X1 OAI21X1_3926 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_0_), .B(_9247_), .C(_9248_), .Y(_9249_) );
	NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_csr_wr), .B(csr_gpr_iu_csr_ret), .Y(_9250_) );
	NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_9250_), .B(_6759__bF_buf3), .Y(_9251_) );
	OAI21X1 OAI21X1_3927 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_9149__bF_buf2), .C(_9251__bF_buf6), .Y(_9252_) );
	OAI21X1 OAI21X1_3928 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_0_), .B(_9251__bF_buf5), .C(_9252_), .Y(_9253_) );
	AOI22X1 AOI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .B(_9097_), .C(csr_gpr_iu_csr_sepc_0_), .D(_9098__bF_buf2), .Y(_9254_) );
	OAI21X1 OAI21X1_3929 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_9105__bF_buf2), .C(_9254_), .Y(_9255_) );
	NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_9094__bF_buf0), .Y(_9256_) );
	OAI21X1 OAI21X1_3930 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf5), .B(_9253_), .C(_9256_), .Y(_9257_) );
	OAI21X1 OAI21X1_3931 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf10_bF_buf1), .B(_9257_), .C(_6879__bF_buf16), .Y(_9258_) );
	AOI21X1 AOI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_9249_), .B(_7303__bF_buf9_bF_buf1), .C(_9258_), .Y(_6725__0_) );
	NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_9247_), .Y(_9259_) );
	OAI21X1 OAI21X1_3932 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_1_), .B(_9247_), .C(_9259_), .Y(_9260_) );
	OAI21X1 OAI21X1_3933 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_9149__bF_buf1), .C(_9251__bF_buf4), .Y(_9261_) );
	OAI21X1 OAI21X1_3934 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_1_), .B(_9251__bF_buf3), .C(_9261_), .Y(_9262_) );
	AOI22X1 AOI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .B(_9097_), .C(csr_gpr_iu_csr_sepc_1_), .D(_9098__bF_buf1), .Y(_9263_) );
	OAI21X1 OAI21X1_3935 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .B(_9105__bF_buf1), .C(_9263_), .Y(_9264_) );
	NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_9264_), .B(_9094__bF_buf4), .Y(_9265_) );
	OAI21X1 OAI21X1_3936 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf3), .B(_9262_), .C(_9265_), .Y(_9266_) );
	OAI21X1 OAI21X1_3937 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf8_bF_buf1), .B(_9266_), .C(_6879__bF_buf15), .Y(_9267_) );
	AOI21X1 AOI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_7303__bF_buf7_bF_buf1), .C(_9267_), .Y(_6725__1_) );
	INVX8 INVX8_85 ( .gnd(gnd), .vdd(vdd), .A(_9247_), .Y(_9268_) );
	INVX1 INVX1_1593 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_2_), .Y(_9269_) );
	AOI21X1 AOI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf6), .B(_9269_), .C(_7304__bF_buf1), .Y(_9270_) );
	OAI21X1 OAI21X1_3938 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(_9268__bF_buf5), .C(_9270_), .Y(_9271_) );
	INVX1 INVX1_1594 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_2_), .Y(_9272_) );
	NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_0_), .B(csr_gpr_iu_csr_mtvec_1_), .Y(_9273_) );
	INVX4 INVX4_21 ( .gnd(gnd), .vdd(vdd), .A(_9273__bF_buf3), .Y(_9274_) );
	OAI21X1 OAI21X1_3939 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_0_), .B(csr_gpr_iu_csr_mtvec_1_), .C(csr_gpr_iu_csr_mcause_31_), .Y(_9275_) );
	INVX4 INVX4_22 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .Y(_9276_) );
	OAI21X1 OAI21X1_3940 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_9272_), .C(_9276__bF_buf3), .Y(_9277_) );
	OAI21X1 OAI21X1_3941 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(_9274_), .C(_9277_), .Y(_9278_) );
	OAI21X1 OAI21X1_3942 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_0_), .B(csr_gpr_iu_csr_mtvec_2_), .C(_9278_), .Y(_9279_) );
	OAI21X1 OAI21X1_3943 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_0_), .B(csr_gpr_iu_csr_mtvec_1_), .C(_8840_), .Y(_9280_) );
	INVX8 INVX8_86 ( .gnd(gnd), .vdd(vdd), .A(_9280_), .Y(_9281_) );
	AOI21X1 AOI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_3_), .B(_9281__bF_buf3), .C(_8861__bF_buf0), .Y(_9282_) );
	INVX1 INVX1_1595 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_2_), .Y(_9283_) );
	NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_0_), .B(csr_gpr_iu_csr_stvec_1_), .Y(_9284_) );
	INVX8 INVX8_87 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .Y(_9285_) );
	NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_9283_), .Y(_9286_) );
	NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_0_), .B(csr_gpr_iu_csr_stvec_2_), .Y(_9287_) );
	AOI21X1 AOI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_9287_), .C(_7571_), .Y(_9288_) );
	OAI21X1 OAI21X1_3944 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf2), .B(csr_gpr_iu_csr_stvec_3_), .C(_9285__bF_buf4), .Y(_9289_) );
	OAI22X1 OAI22X1_746 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .B(_9285__bF_buf3), .C(_9289_), .D(_9288_), .Y(_9290_) );
	INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(_9149__bF_buf0), .Y(_9291_) );
	INVX4 INVX4_23 ( .gnd(gnd), .vdd(vdd), .A(_9251__bF_buf2), .Y(_9292_) );
	AOI21X1 AOI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_7595_), .C(_9292_), .Y(_9293_) );
	OAI21X1 OAI21X1_3945 ( .gnd(gnd), .vdd(vdd), .A(_7594__bF_buf5), .B(_9290_), .C(_9293_), .Y(_9294_) );
	AOI21X1 AOI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_9279_), .B(_9282_), .C(_9294_), .Y(_9295_) );
	OAI21X1 OAI21X1_3946 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(_9251__bF_buf1), .C(_9095__bF_buf0), .Y(_9296_) );
	AOI22X1 AOI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(_9097_), .C(csr_gpr_iu_csr_sepc_2_), .D(_9098__bF_buf0), .Y(_9297_) );
	OAI21X1 OAI21X1_3947 ( .gnd(gnd), .vdd(vdd), .A(_8858_), .B(_9105__bF_buf0), .C(_9297_), .Y(_9298_) );
	INVX1 INVX1_1596 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9299_) );
	AOI21X1 AOI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf2), .B(_9299_), .C(_7303__bF_buf6_bF_buf1), .Y(_9300_) );
	OAI21X1 OAI21X1_3948 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_9295_), .C(_9300_), .Y(_9301_) );
	AOI21X1 AOI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_9271_), .B(_9301_), .C(rst_bF_buf44), .Y(_6725__2_) );
	INVX1 INVX1_1597 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_3_), .Y(_9302_) );
	AOI21X1 AOI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf4), .B(_9302_), .C(_7304__bF_buf0), .Y(_9303_) );
	OAI21X1 OAI21X1_3949 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .B(_9268__bF_buf3), .C(_9303_), .Y(_9304_) );
	NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_0_), .B(csr_gpr_iu_csr_mtvec_2_), .Y(_9305_) );
	NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .B(csr_gpr_iu_csr_mtvec_3_), .Y(_9306_) );
	INVX1 INVX1_1598 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9307_) );
	NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .B(csr_gpr_iu_csr_mtvec_3_), .Y(_9308_) );
	NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_9307_), .Y(_9309_) );
	NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .B(_9309_), .Y(_9310_) );
	OAI21X1 OAI21X1_3950 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_9272_), .C(_9309_), .Y(_9311_) );
	NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf2), .B(_9311_), .Y(_9312_) );
	AOI22X1 AOI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_3_), .B(_9273__bF_buf2), .C(csr_gpr_iu_csr_mtvec_4_), .D(_9281__bF_buf2), .Y(_9313_) );
	OAI21X1 OAI21X1_3951 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .B(_9312_), .C(_9313_), .Y(_9314_) );
	INVX1 INVX1_1599 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9315_) );
	NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .B(csr_gpr_iu_csr_stvec_3_), .Y(_9316_) );
	NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_1_), .B(csr_gpr_iu_csr_stvec_3_), .Y(_9317_) );
	INVX1 INVX1_1600 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9318_) );
	NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .B(_9318_), .Y(_9319_) );
	NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_9319_), .Y(_9320_) );
	OAI21X1 OAI21X1_3952 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_0_), .B(csr_gpr_iu_csr_stvec_1_), .C(csr_gpr_iu_csr_scause_31_bF_buf1), .Y(_9321_) );
	INVX4 INVX4_24 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_9322_) );
	INVX1 INVX1_1601 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .Y(_9323_) );
	OAI21X1 OAI21X1_3953 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .B(_9323_), .C(_9322__bF_buf3), .Y(_9324_) );
	OAI21X1 OAI21X1_3954 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_0_), .B(csr_gpr_iu_csr_stvec_1_), .C(_7571_), .Y(_9325_) );
	INVX4 INVX4_25 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9326_) );
	INVX1 INVX1_1602 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_3_), .Y(_9327_) );
	OAI21X1 OAI21X1_3955 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9285__bF_buf2), .C(_9149__bF_buf4), .Y(_9328_) );
	AOI21X1 AOI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_4_), .B(_9326_), .C(_9328_), .Y(_9329_) );
	OAI21X1 OAI21X1_3956 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9324_), .C(_9329_), .Y(_9330_) );
	AOI22X1 AOI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf1), .B(_9314_), .C(_8861__bF_buf6), .D(_9330_), .Y(_9331_) );
	OAI21X1 OAI21X1_3957 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .B(_9149__bF_buf3), .C(_9251__bF_buf0), .Y(_9332_) );
	NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_9332_), .B(_9331_), .Y(_9333_) );
	OAI21X1 OAI21X1_3958 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_9251__bF_buf6), .C(_9095__bF_buf4), .Y(_9334_) );
	AOI22X1 AOI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .B(_9097_), .C(csr_gpr_iu_csr_sepc_3_), .D(_9098__bF_buf4), .Y(_9335_) );
	OAI21X1 OAI21X1_3959 ( .gnd(gnd), .vdd(vdd), .A(_8864_), .B(_9105__bF_buf4), .C(_9335_), .Y(_9336_) );
	INVX1 INVX1_1603 ( .gnd(gnd), .vdd(vdd), .A(_9336_), .Y(_9337_) );
	AOI21X1 AOI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf1), .B(_9337_), .C(_7303__bF_buf5_bF_buf1), .Y(_9338_) );
	OAI21X1 OAI21X1_3960 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .B(_9333_), .C(_9338_), .Y(_9339_) );
	AOI21X1 AOI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_9339_), .C(rst_bF_buf43), .Y(_6725__3_) );
	INVX1 INVX1_1604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_4_), .Y(_9340_) );
	AOI21X1 AOI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf2), .B(_9340_), .C(_7304__bF_buf14_bF_buf0), .Y(_9341_) );
	OAI21X1 OAI21X1_3961 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .B(_9268__bF_buf1), .C(_9341_), .Y(_9342_) );
	OAI21X1 OAI21X1_3962 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .B(_9306_), .C(_9308_), .Y(_9343_) );
	INVX1 INVX1_1605 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_4_), .Y(_9344_) );
	NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_9344_), .Y(_9345_) );
	NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .B(csr_gpr_iu_csr_mtvec_4_), .Y(_9346_) );
	NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_9346_), .B(_9345_), .Y(_9347_) );
	INVX1 INVX1_1606 ( .gnd(gnd), .vdd(vdd), .A(_9347_), .Y(_9348_) );
	AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_9348_), .B(_9343_), .Y(_9349_) );
	OAI21X1 OAI21X1_3963 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9348_), .C(_9276__bF_buf1), .Y(_9350_) );
	AOI22X1 AOI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_4_), .B(_9273__bF_buf1), .C(csr_gpr_iu_csr_mtvec_5_), .D(_9281__bF_buf1), .Y(_9351_) );
	OAI21X1 OAI21X1_3964 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_9350_), .C(_9351_), .Y(_9352_) );
	OAI21X1 OAI21X1_3965 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .B(_9316_), .C(_9317_), .Y(_9353_) );
	NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .B(csr_gpr_iu_csr_stvec_4_), .Y(_9354_) );
	AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .B(csr_gpr_iu_csr_stvec_4_), .Y(_9355_) );
	NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_9355_), .Y(_9356_) );
	NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9353_), .Y(_9357_) );
	NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9353_), .Y(_9358_) );
	NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf2), .B(_9358_), .Y(_9359_) );
	INVX1 INVX1_1607 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_4_), .Y(_9360_) );
	OAI21X1 OAI21X1_3966 ( .gnd(gnd), .vdd(vdd), .A(_9360_), .B(_9285__bF_buf1), .C(_9149__bF_buf2), .Y(_9361_) );
	AOI21X1 AOI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_5_), .B(_9326_), .C(_9361_), .Y(_9362_) );
	OAI21X1 OAI21X1_3967 ( .gnd(gnd), .vdd(vdd), .A(_9357_), .B(_9359_), .C(_9362_), .Y(_9363_) );
	AOI22X1 AOI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf0), .B(_9352_), .C(_8861__bF_buf5), .D(_9363_), .Y(_9364_) );
	OAI21X1 OAI21X1_3968 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .B(_9149__bF_buf1), .C(_9251__bF_buf5), .Y(_9365_) );
	NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_9364_), .Y(_9366_) );
	OAI21X1 OAI21X1_3969 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_9251__bF_buf4), .C(_9095__bF_buf3), .Y(_9367_) );
	OAI22X1 OAI22X1_747 ( .gnd(gnd), .vdd(vdd), .A(_7645_), .B(biu_mmu_msu_0_bF_buf1), .C(_8869_), .D(_9105__bF_buf3), .Y(_9368_) );
	AOI21X1 AOI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_4_), .B(_9098__bF_buf3), .C(_9368_), .Y(_9369_) );
	AOI21X1 AOI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_9369_), .B(_9094__bF_buf0), .C(_7303__bF_buf4_bF_buf1), .Y(_9370_) );
	OAI21X1 OAI21X1_3970 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_9366_), .C(_9370_), .Y(_9371_) );
	AOI21X1 AOI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9371_), .C(rst_bF_buf42), .Y(_6725__4_) );
	INVX1 INVX1_1608 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_5_), .Y(_9372_) );
	AOI21X1 AOI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf0), .B(_9372_), .C(_7304__bF_buf13_bF_buf0), .Y(_9373_) );
	OAI21X1 OAI21X1_3971 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .B(_9268__bF_buf6), .C(_9373_), .Y(_9374_) );
	OAI21X1 OAI21X1_3972 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf0), .B(csr_gpr_iu_csr_stvec_6_), .C(_9285__bF_buf0), .Y(_9375_) );
	OAI21X1 OAI21X1_3973 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_9360_), .C(_9358_), .Y(_9376_) );
	NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_3_), .B(csr_gpr_iu_csr_stvec_5_), .Y(_9377_) );
	AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_3_), .B(csr_gpr_iu_csr_stvec_5_), .Y(_9378_) );
	NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_9377_), .B(_9378_), .Y(_9379_) );
	XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_9379_), .Y(_9380_) );
	AOI21X1 AOI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_9380_), .B(csr_gpr_iu_csr_scause_31_bF_buf3), .C(_9375_), .Y(_9381_) );
	INVX1 INVX1_1609 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_5_), .Y(_9382_) );
	OAI21X1 OAI21X1_3974 ( .gnd(gnd), .vdd(vdd), .A(_9382_), .B(_9285__bF_buf4), .C(_9149__bF_buf0), .Y(_9383_) );
	OAI21X1 OAI21X1_3975 ( .gnd(gnd), .vdd(vdd), .A(_9383_), .B(_9381_), .C(_8861__bF_buf4), .Y(_9384_) );
	INVX1 INVX1_1610 ( .gnd(gnd), .vdd(vdd), .A(_9346_), .Y(_9385_) );
	NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_9385_), .B(_9349_), .Y(_9386_) );
	INVX1 INVX1_1611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_5_), .Y(_9387_) );
	NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_9387_), .Y(_9388_) );
	NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_3_), .B(csr_gpr_iu_csr_mtvec_5_), .Y(_9389_) );
	NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_9389_), .B(_9388_), .Y(_9390_) );
	NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_9386_), .Y(_9391_) );
	INVX1 INVX1_1612 ( .gnd(gnd), .vdd(vdd), .A(_9386_), .Y(_9392_) );
	INVX1 INVX1_1613 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .Y(_9393_) );
	OAI21X1 OAI21X1_3976 ( .gnd(gnd), .vdd(vdd), .A(_9393_), .B(_9392_), .C(_9276__bF_buf0), .Y(_9394_) );
	AOI22X1 AOI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_5_), .B(_9273__bF_buf0), .C(csr_gpr_iu_csr_mtvec_6_), .D(_9281__bF_buf0), .Y(_9395_) );
	OAI21X1 OAI21X1_3977 ( .gnd(gnd), .vdd(vdd), .A(_9391_), .B(_9394_), .C(_9395_), .Y(_9396_) );
	NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf3), .B(_9396_), .Y(_9397_) );
	OAI21X1 OAI21X1_3978 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .B(_9149__bF_buf4), .C(_9251__bF_buf3), .Y(_9398_) );
	AOI21X1 AOI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_9397_), .B(_9384_), .C(_9398_), .Y(_9399_) );
	OAI21X1 OAI21X1_3979 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .B(_9251__bF_buf2), .C(_9095__bF_buf2), .Y(_9400_) );
	OAI22X1 OAI22X1_748 ( .gnd(gnd), .vdd(vdd), .A(_7656_), .B(biu_mmu_msu_0_bF_buf0), .C(_8874_), .D(_9105__bF_buf2), .Y(_9401_) );
	AOI21X1 AOI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_5_), .B(_9098__bF_buf2), .C(_9401_), .Y(_9402_) );
	AOI21X1 AOI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_9402_), .B(_9094__bF_buf5), .C(_7303__bF_buf3_bF_buf1), .Y(_9403_) );
	OAI21X1 OAI21X1_3980 ( .gnd(gnd), .vdd(vdd), .A(_9400_), .B(_9399_), .C(_9403_), .Y(_9404_) );
	AOI21X1 AOI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .B(_9404_), .C(rst_bF_buf41), .Y(_6725__5_) );
	AOI22X1 AOI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .B(_9097_), .C(csr_gpr_iu_csr_sepc_6_), .D(_9098__bF_buf1), .Y(_9405_) );
	OAI21X1 OAI21X1_3981 ( .gnd(gnd), .vdd(vdd), .A(_8882_), .B(_9105__bF_buf1), .C(_9405_), .Y(_9406_) );
	INVX1 INVX1_1614 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_6_), .Y(_9407_) );
	OAI21X1 OAI21X1_3982 ( .gnd(gnd), .vdd(vdd), .A(_9407_), .B(_9285__bF_buf3), .C(_9149__bF_buf3), .Y(_9408_) );
	NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .B(csr_gpr_iu_csr_stvec_6_), .Y(_9409_) );
	AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .B(csr_gpr_iu_csr_stvec_6_), .Y(_9410_) );
	NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_9409_), .B(_9410_), .Y(_9411_) );
	NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9353_), .C(_9379_), .Y(_9412_) );
	NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .B(csr_gpr_iu_csr_stvec_4_), .Y(_9413_) );
	NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_3_), .B(csr_gpr_iu_csr_stvec_5_), .Y(_9414_) );
	OAI21X1 OAI21X1_3983 ( .gnd(gnd), .vdd(vdd), .A(_9413_), .B(_9377_), .C(_9414_), .Y(_9415_) );
	INVX1 INVX1_1615 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .Y(_9416_) );
	NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_9416_), .B(_9412_), .Y(_9417_) );
	XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_9417_), .B(_9411_), .Y(_9418_) );
	OAI21X1 OAI21X1_3984 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf2), .B(csr_gpr_iu_csr_stvec_7_), .C(_9285__bF_buf2), .Y(_9419_) );
	AOI21X1 AOI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_9418_), .B(csr_gpr_iu_csr_scause_31_bF_buf1), .C(_9419_), .Y(_9420_) );
	OAI21X1 OAI21X1_3985 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .B(_9420_), .C(_8861__bF_buf3), .Y(_9421_) );
	INVX1 INVX1_1616 ( .gnd(gnd), .vdd(vdd), .A(_9388_), .Y(_9422_) );
	OAI21X1 OAI21X1_3986 ( .gnd(gnd), .vdd(vdd), .A(_9346_), .B(_9422_), .C(_9389_), .Y(_9423_) );
	INVX1 INVX1_1617 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .Y(_9424_) );
	NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_9347_), .B(_9390_), .Y(_9425_) );
	NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9425_), .Y(_9426_) );
	NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_9424_), .B(_9426_), .Y(_9427_) );
	INVX1 INVX1_1618 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_6_), .Y(_9428_) );
	NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_9428_), .Y(_9429_) );
	NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .B(csr_gpr_iu_csr_mtvec_6_), .Y(_9430_) );
	NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_9430_), .B(_9429_), .Y(_9431_) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_9427_), .B(_9431_), .Y(_9432_) );
	AOI22X1 AOI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_6_), .B(_9273__bF_buf3), .C(csr_gpr_iu_csr_mtvec_7_), .D(_9281__bF_buf3), .Y(_9433_) );
	OAI21X1 OAI21X1_3987 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_9432_), .C(_9433_), .Y(_9434_) );
	NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf2), .B(_9434_), .Y(_9435_) );
	OAI21X1 OAI21X1_3988 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .B(_9149__bF_buf2), .C(_9251__bF_buf1), .Y(_9436_) );
	AOI21X1 AOI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_9435_), .B(_9421_), .C(_9436_), .Y(_9437_) );
	INVX1 INVX1_1619 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_6_), .Y(_9438_) );
	OAI21X1 OAI21X1_3989 ( .gnd(gnd), .vdd(vdd), .A(_9438_), .B(_9251__bF_buf0), .C(_9095__bF_buf1), .Y(_9439_) );
	OAI22X1 OAI22X1_749 ( .gnd(gnd), .vdd(vdd), .A(_9095__bF_buf0), .B(_9406_), .C(_9439_), .D(_9437_), .Y(_9440_) );
	NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_7666_), .B(_9268__bF_buf5), .Y(_9441_) );
	OAI21X1 OAI21X1_3990 ( .gnd(gnd), .vdd(vdd), .A(_9438_), .B(_9247_), .C(_7303__bF_buf2), .Y(_9442_) );
	OAI21X1 OAI21X1_3991 ( .gnd(gnd), .vdd(vdd), .A(_9442_), .B(_9441_), .C(_6879__bF_buf14), .Y(_9443_) );
	AOI21X1 AOI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_9440_), .B(_7304__bF_buf12_bF_buf0), .C(_9443_), .Y(_6725__6_) );
	INVX1 INVX1_1620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_7_), .Y(_9444_) );
	AOI21X1 AOI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf4), .B(_9444_), .C(_7304__bF_buf11_bF_buf0), .Y(_9445_) );
	OAI21X1 OAI21X1_3992 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .B(_9268__bF_buf3), .C(_9445_), .Y(_9446_) );
	OAI21X1 OAI21X1_3993 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf0), .B(csr_gpr_iu_csr_stvec_8_), .C(_9285__bF_buf1), .Y(_9447_) );
	AOI21X1 AOI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_9417_), .B(_9411_), .C(_9410_), .Y(_9448_) );
	NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .B(csr_gpr_iu_csr_stvec_7_), .Y(_9449_) );
	AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .B(csr_gpr_iu_csr_stvec_7_), .Y(_9450_) );
	NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_9449_), .B(_9450_), .Y(_9451_) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_9448_), .B(_9451_), .Y(_9452_) );
	AOI21X1 AOI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_9452_), .B(csr_gpr_iu_csr_scause_31_bF_buf3), .C(_9447_), .Y(_9453_) );
	INVX1 INVX1_1621 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_7_), .Y(_9454_) );
	OAI21X1 OAI21X1_3994 ( .gnd(gnd), .vdd(vdd), .A(_9454_), .B(_9285__bF_buf0), .C(_7426_), .Y(_9455_) );
	AOI21X1 AOI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7673_), .C(_8614_), .Y(_9456_) );
	OAI21X1 OAI21X1_3995 ( .gnd(gnd), .vdd(vdd), .A(_9455_), .B(_9453_), .C(_9456_), .Y(_9457_) );
	INVX1 INVX1_1622 ( .gnd(gnd), .vdd(vdd), .A(_9427_), .Y(_9458_) );
	OAI21X1 OAI21X1_3996 ( .gnd(gnd), .vdd(vdd), .A(_9431_), .B(_9458_), .C(_9430_), .Y(_9459_) );
	OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .B(csr_gpr_iu_csr_mtvec_7_), .Y(_9460_) );
	NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf5), .B(csr_gpr_iu_csr_mtvec_7_), .Y(_9461_) );
	NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_9461_), .B(_9460_), .Y(_9462_) );
	XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9462_), .Y(_9463_) );
	AOI22X1 AOI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_7_), .B(_9273__bF_buf2), .C(csr_gpr_iu_csr_mtvec_8_), .D(_9281__bF_buf2), .Y(_9464_) );
	OAI21X1 OAI21X1_3997 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_9463_), .C(_9464_), .Y(_9465_) );
	AOI21X1 AOI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_8614_), .C(_7424__bF_buf0), .Y(_9466_) );
	OAI21X1 OAI21X1_3998 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .B(_7423_), .C(_9251__bF_buf6), .Y(_9467_) );
	AOI21X1 AOI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_9457_), .C(_9467_), .Y(_9468_) );
	OAI21X1 OAI21X1_3999 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_9251__bF_buf5), .C(_9095__bF_buf4), .Y(_9469_) );
	OAI22X1 OAI22X1_750 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(biu_mmu_msu_0_bF_buf4), .C(_8885_), .D(_9105__bF_buf0), .Y(_9470_) );
	AOI21X1 AOI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_7_), .B(_9098__bF_buf0), .C(_9470_), .Y(_9471_) );
	AOI21X1 AOI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_9471_), .B(_9094__bF_buf4), .C(_7303__bF_buf1), .Y(_9472_) );
	OAI21X1 OAI21X1_4000 ( .gnd(gnd), .vdd(vdd), .A(_9469_), .B(_9468_), .C(_9472_), .Y(_9473_) );
	AOI21X1 AOI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_9473_), .B(_9446_), .C(rst_bF_buf40), .Y(_6725__7_) );
	INVX1 INVX1_1623 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_8_), .Y(_9474_) );
	AOI21X1 AOI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf2), .B(_9474_), .C(_7304__bF_buf10_bF_buf0), .Y(_9475_) );
	OAI21X1 OAI21X1_4001 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .B(_9268__bF_buf1), .C(_9475_), .Y(_9476_) );
	INVX1 INVX1_1624 ( .gnd(gnd), .vdd(vdd), .A(_9449_), .Y(_9477_) );
	AOI21X1 AOI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_9477_), .B(_9410_), .C(_9450_), .Y(_9478_) );
	NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9415_), .C(_9451_), .Y(_9479_) );
	AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_9479_), .B(_9478_), .Y(_9480_) );
	OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_2_), .B(csr_gpr_iu_csr_stvec_4_), .Y(_9481_) );
	NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_9413_), .B(_9481_), .Y(_9482_) );
	NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_9382_), .Y(_9483_) );
	NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_9414_), .B(_9483_), .Y(_9484_) );
	NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_9484_), .Y(_9485_) );
	AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9451_), .Y(_9486_) );
	NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_9485_), .C(_9486_), .Y(_9487_) );
	NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_9487_), .B(_9480_), .Y(_9488_) );
	OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf4), .B(csr_gpr_iu_csr_stvec_8_), .Y(_9489_) );
	NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf3), .B(csr_gpr_iu_csr_stvec_8_), .Y(_9490_) );
	NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_9490_), .B(_9489_), .Y(_9491_) );
	INVX1 INVX1_1625 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .Y(_9492_) );
	OAI21X1 OAI21X1_4002 ( .gnd(gnd), .vdd(vdd), .A(_9492_), .B(_9488_), .C(_9322__bF_buf1), .Y(_9493_) );
	AOI21X1 AOI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .B(_9492_), .C(_9493_), .Y(_9494_) );
	INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_9_), .Y(_9495_) );
	AOI21X1 AOI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_8_), .B(_9284_), .C(_9291_), .Y(_9496_) );
	OAI21X1 OAI21X1_4003 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9325_), .C(_9496_), .Y(_9497_) );
	OAI21X1 OAI21X1_4004 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_9494_), .C(_8861__bF_buf2), .Y(_9498_) );
	OAI21X1 OAI21X1_4005 ( .gnd(gnd), .vdd(vdd), .A(_9430_), .B(_9462_), .C(_9461_), .Y(_9499_) );
	NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_9462_), .B(_9431_), .Y(_9500_) );
	AOI21X1 AOI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_9500_), .C(_9499_), .Y(_9501_) );
	NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9500_), .C(_9425_), .Y(_9502_) );
	NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_9502_), .B(_9501_), .Y(_9503_) );
	INVX1 INVX1_1626 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .Y(_9504_) );
	INVX1 INVX1_1627 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_8_), .Y(_9505_) );
	NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_9505_), .Y(_9506_) );
	NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf2), .B(csr_gpr_iu_csr_mtvec_8_), .Y(_9507_) );
	NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_9507_), .B(_9506_), .Y(_9508_) );
	NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_9508_), .B(_9504_), .Y(_9509_) );
	INVX1 INVX1_1628 ( .gnd(gnd), .vdd(vdd), .A(_9508_), .Y(_9510_) );
	OAI21X1 OAI21X1_4006 ( .gnd(gnd), .vdd(vdd), .A(_9510_), .B(_9503_), .C(_9276__bF_buf3), .Y(_9511_) );
	AOI22X1 AOI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_8_), .B(_9273__bF_buf1), .C(csr_gpr_iu_csr_mtvec_9_), .D(_9281__bF_buf1), .Y(_9512_) );
	OAI21X1 OAI21X1_4007 ( .gnd(gnd), .vdd(vdd), .A(_9511_), .B(_9509_), .C(_9512_), .Y(_9513_) );
	NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf1), .B(_9513_), .Y(_9514_) );
	OAI21X1 OAI21X1_4008 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .B(_9149__bF_buf1), .C(_9251__bF_buf4), .Y(_9515_) );
	AOI21X1 AOI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_9514_), .B(_9498_), .C(_9515_), .Y(_9516_) );
	OAI21X1 OAI21X1_4009 ( .gnd(gnd), .vdd(vdd), .A(_9474_), .B(_9251__bF_buf3), .C(_9095__bF_buf3), .Y(_9517_) );
	OAI22X1 OAI22X1_751 ( .gnd(gnd), .vdd(vdd), .A(_7699_), .B(biu_mmu_msu_0_bF_buf3), .C(_8890_), .D(_9105__bF_buf4), .Y(_9518_) );
	AOI21X1 AOI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_8_), .B(_9098__bF_buf4), .C(_9518_), .Y(_9519_) );
	AOI21X1 AOI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_9519_), .B(_9094__bF_buf3), .C(_7303__bF_buf0), .Y(_9520_) );
	OAI21X1 OAI21X1_4010 ( .gnd(gnd), .vdd(vdd), .A(_9517_), .B(_9516_), .C(_9520_), .Y(_9521_) );
	AOI21X1 AOI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_9476_), .B(_9521_), .C(rst_bF_buf39), .Y(_6725__8_) );
	INVX1 INVX1_1629 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_9_), .Y(_9522_) );
	AOI21X1 AOI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf0), .B(_9522_), .C(_7304__bF_buf9_bF_buf0), .Y(_9523_) );
	OAI21X1 OAI21X1_4011 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .B(_9268__bF_buf6), .C(_9523_), .Y(_9524_) );
	OAI21X1 OAI21X1_4012 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf2), .B(csr_gpr_iu_csr_stvec_10_), .C(_9285__bF_buf4), .Y(_9525_) );
	INVX1 INVX1_1630 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .Y(_9526_) );
	AOI21X1 AOI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_9417_), .B(_9486_), .C(_9526_), .Y(_9527_) );
	OAI21X1 OAI21X1_4013 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(_9527_), .C(_9490_), .Y(_9528_) );
	NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .B(_9495_), .Y(_9529_) );
	NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf1), .B(csr_gpr_iu_csr_stvec_9_), .Y(_9530_) );
	NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_9530_), .B(_9529_), .Y(_9531_) );
	INVX1 INVX1_1631 ( .gnd(gnd), .vdd(vdd), .A(_9531_), .Y(_9532_) );
	XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_9528_), .B(_9532_), .Y(_9533_) );
	AOI21X1 AOI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(csr_gpr_iu_csr_scause_31_bF_buf1), .C(_9525_), .Y(_9534_) );
	OAI21X1 OAI21X1_4014 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9285__bF_buf3), .C(_9149__bF_buf0), .Y(_9535_) );
	OAI21X1 OAI21X1_4015 ( .gnd(gnd), .vdd(vdd), .A(_9535_), .B(_9534_), .C(_8861__bF_buf1), .Y(_9536_) );
	AOI21X1 AOI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf0), .B(csr_gpr_iu_csr_mtvec_8_), .C(_9509_), .Y(_9537_) );
	INVX1 INVX1_1632 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_9_), .Y(_9538_) );
	NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .B(_9538_), .Y(_9539_) );
	NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_cause_31_bF_buf6), .B(csr_gpr_iu_csr_mtvec_9_), .Y(_9540_) );
	NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9539_), .Y(_9541_) );
	INVX1 INVX1_1633 ( .gnd(gnd), .vdd(vdd), .A(_9541_), .Y(_9542_) );
	AOI21X1 AOI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_9537_), .B(_9542_), .C(_9275_), .Y(_9543_) );
	OAI21X1 OAI21X1_4016 ( .gnd(gnd), .vdd(vdd), .A(_9537_), .B(_9542_), .C(_9543_), .Y(_9544_) );
	INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_10_), .Y(_9545_) );
	OAI21X1 OAI21X1_4017 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_9_), .B(_9274_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf0), .Y(_9546_) );
	AOI21X1 AOI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_9545_), .B(_9281__bF_buf0), .C(_9546_), .Y(_9547_) );
	NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_9547_), .B(_9544_), .Y(_9548_) );
	OAI21X1 OAI21X1_4018 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .B(_9149__bF_buf4), .C(_9251__bF_buf2), .Y(_9549_) );
	AOI21X1 AOI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_9548_), .B(_9536_), .C(_9549_), .Y(_9550_) );
	OAI21X1 OAI21X1_4019 ( .gnd(gnd), .vdd(vdd), .A(_9522_), .B(_9251__bF_buf1), .C(_9095__bF_buf2), .Y(_9551_) );
	OAI22X1 OAI22X1_752 ( .gnd(gnd), .vdd(vdd), .A(_7698_), .B(biu_mmu_msu_0_bF_buf2), .C(_8897_), .D(_9105__bF_buf3), .Y(_9552_) );
	AOI21X1 AOI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_9_), .B(_9098__bF_buf3), .C(_9552_), .Y(_9553_) );
	AOI21X1 AOI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_9553_), .B(_9094__bF_buf2), .C(_7303__bF_buf14_bF_buf0), .Y(_9554_) );
	OAI21X1 OAI21X1_4020 ( .gnd(gnd), .vdd(vdd), .A(_9551_), .B(_9550_), .C(_9554_), .Y(_9555_) );
	AOI21X1 AOI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_9555_), .B(_9524_), .C(rst_bF_buf38), .Y(_6725__9_) );
	INVX1 INVX1_1634 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_10_), .Y(_9556_) );
	AOI21X1 AOI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf5), .B(_9556_), .C(_7304__bF_buf8_bF_buf0), .Y(_9557_) );
	OAI21X1 OAI21X1_4021 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(_9268__bF_buf4), .C(_9557_), .Y(_9558_) );
	OAI21X1 OAI21X1_4022 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7709_), .C(_7427_), .Y(_9559_) );
	NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(_9531_), .Y(_9560_) );
	INVX1 INVX1_1635 ( .gnd(gnd), .vdd(vdd), .A(_9560_), .Y(_9561_) );
	OAI21X1 OAI21X1_4023 ( .gnd(gnd), .vdd(vdd), .A(_9490_), .B(_9531_), .C(_9530_), .Y(_9562_) );
	INVX1 INVX1_1636 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .Y(_9563_) );
	OAI21X1 OAI21X1_4024 ( .gnd(gnd), .vdd(vdd), .A(_9561_), .B(_9527_), .C(_9563_), .Y(_9564_) );
	OAI21X1 OAI21X1_4025 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_10_), .B(_9564_), .C(_9322__bF_buf0), .Y(_9565_) );
	AOI21X1 AOI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_10_), .B(_9564_), .C(_9565_), .Y(_9566_) );
	INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_11_), .Y(_9567_) );
	AOI21X1 AOI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_10_), .B(_9284_), .C(_7427_), .Y(_9568_) );
	OAI21X1 OAI21X1_4026 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_9325_), .C(_9568_), .Y(_9569_) );
	OAI21X1 OAI21X1_4027 ( .gnd(gnd), .vdd(vdd), .A(_9569_), .B(_9566_), .C(_9559_), .Y(_9570_) );
	NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_9508_), .B(_9541_), .Y(_9571_) );
	OAI21X1 OAI21X1_4028 ( .gnd(gnd), .vdd(vdd), .A(_9507_), .B(_9541_), .C(_9540_), .Y(_9572_) );
	AOI21X1 AOI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .B(_9571_), .C(_9572_), .Y(_9573_) );
	NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_9545_), .B(_9573_), .Y(_9574_) );
	NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_9545_), .B(_9573_), .Y(_9575_) );
	INVX1 INVX1_1637 ( .gnd(gnd), .vdd(vdd), .A(_9575_), .Y(_9576_) );
	NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_9574_), .B(_9576_), .Y(_9577_) );
	AOI22X1 AOI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_10_), .B(_9273__bF_buf0), .C(csr_gpr_iu_csr_mtvec_11_), .D(_9281__bF_buf3), .Y(_9578_) );
	OAI21X1 OAI21X1_4029 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_9577_), .C(_9578_), .Y(_9579_) );
	AOI21X1 AOI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_9579_), .B(_8614_), .C(_7424__bF_buf3), .Y(_9580_) );
	OAI21X1 OAI21X1_4030 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(_7423_), .C(_9251__bF_buf0), .Y(_9581_) );
	AOI21X1 AOI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_9580_), .B(_9570_), .C(_9581_), .Y(_9582_) );
	OAI21X1 OAI21X1_4031 ( .gnd(gnd), .vdd(vdd), .A(_9556_), .B(_9251__bF_buf6), .C(_9095__bF_buf1), .Y(_9583_) );
	OAI22X1 OAI22X1_753 ( .gnd(gnd), .vdd(vdd), .A(_7709_), .B(biu_mmu_msu_0_bF_buf1), .C(_8902_), .D(_9105__bF_buf2), .Y(_9584_) );
	AOI21X1 AOI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_10_), .B(_9098__bF_buf2), .C(_9584_), .Y(_9585_) );
	AOI21X1 AOI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_9585_), .B(_9094__bF_buf1), .C(_7303__bF_buf13_bF_buf0), .Y(_9586_) );
	OAI21X1 OAI21X1_4032 ( .gnd(gnd), .vdd(vdd), .A(_9583_), .B(_9582_), .C(_9586_), .Y(_9587_) );
	AOI21X1 AOI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_9587_), .B(_9558_), .C(rst_bF_buf37), .Y(_6725__10_) );
	INVX1 INVX1_1638 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_11_), .Y(_9588_) );
	AOI21X1 AOI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf3), .B(_9588_), .C(_7304__bF_buf7_bF_buf0), .Y(_9589_) );
	OAI21X1 OAI21X1_4033 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(_9268__bF_buf2), .C(_9589_), .Y(_9590_) );
	OAI21X1 OAI21X1_4034 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7723_), .C(_7427_), .Y(_9591_) );
	NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_10_), .B(_9564_), .Y(_9592_) );
	OAI21X1 OAI21X1_4035 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_9592_), .C(_9322__bF_buf3), .Y(_9593_) );
	AOI21X1 AOI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_9592_), .C(_9593_), .Y(_9594_) );
	INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_12_), .Y(_9595_) );
	AOI21X1 AOI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_11_), .B(_9284_), .C(_7427_), .Y(_9596_) );
	OAI21X1 OAI21X1_4036 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9325_), .C(_9596_), .Y(_9597_) );
	OAI21X1 OAI21X1_4037 ( .gnd(gnd), .vdd(vdd), .A(_9597_), .B(_9594_), .C(_9591_), .Y(_9598_) );
	NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_11_), .B(_9575_), .Y(_9599_) );
	INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_11_), .Y(_9600_) );
	OAI21X1 OAI21X1_4038 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_9576_), .C(_9276__bF_buf2), .Y(_9601_) );
	AOI22X1 AOI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_11_), .B(_9273__bF_buf3), .C(csr_gpr_iu_csr_mtvec_12_), .D(_9281__bF_buf2), .Y(_9602_) );
	OAI21X1 OAI21X1_4039 ( .gnd(gnd), .vdd(vdd), .A(_9599_), .B(_9601_), .C(_9602_), .Y(_9603_) );
	AOI21X1 AOI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_9603_), .B(_8614_), .C(_7424__bF_buf2), .Y(_9604_) );
	OAI21X1 OAI21X1_4040 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(_7423_), .C(_9251__bF_buf5), .Y(_9605_) );
	AOI21X1 AOI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_9604_), .B(_9598_), .C(_9605_), .Y(_9606_) );
	OAI21X1 OAI21X1_4041 ( .gnd(gnd), .vdd(vdd), .A(_9588_), .B(_9251__bF_buf4), .C(_9095__bF_buf0), .Y(_9607_) );
	OAI22X1 OAI22X1_754 ( .gnd(gnd), .vdd(vdd), .A(_7723_), .B(biu_mmu_msu_0_bF_buf0), .C(_8907_), .D(_9105__bF_buf1), .Y(_9608_) );
	AOI21X1 AOI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_11_), .B(_9098__bF_buf1), .C(_9608_), .Y(_9609_) );
	AOI21X1 AOI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_9609_), .B(_9094__bF_buf0), .C(_7303__bF_buf12_bF_buf0), .Y(_9610_) );
	OAI21X1 OAI21X1_4042 ( .gnd(gnd), .vdd(vdd), .A(_9607_), .B(_9606_), .C(_9610_), .Y(_9611_) );
	AOI21X1 AOI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_9611_), .B(_9590_), .C(rst_bF_buf36), .Y(_6725__11_) );
	OAI21X1 OAI21X1_4043 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9246_), .C(csr_gpr_iu_csr_pc_next_12_), .Y(_9612_) );
	OAI21X1 OAI21X1_4044 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(_9268__bF_buf1), .C(_9612_), .Y(_9613_) );
	NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf11_bF_buf0), .B(_9613_), .Y(_9614_) );
	INVX1 INVX1_1639 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_12_), .Y(_9615_) );
	OAI21X1 OAI21X1_4045 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_9576_), .C(_9615_), .Y(_9616_) );
	AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_9575_), .B(csr_gpr_iu_csr_mtvec_11_), .Y(_9617_) );
	NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_12_), .B(_9617_), .Y(_9618_) );
	NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf1), .B(_9616_), .C(_9618_), .Y(_9619_) );
	AOI22X1 AOI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_12_), .B(_9273__bF_buf2), .C(csr_gpr_iu_csr_mtvec_13_), .D(_9281__bF_buf1), .Y(_9620_) );
	NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_9620_), .B(_9619_), .Y(_9621_) );
	INVX1 INVX1_1640 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_10_), .Y(_9622_) );
	NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_9622_), .B(_9567_), .Y(_9623_) );
	NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9564_), .Y(_9624_) );
	AOI21X1 AOI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_9624_), .B(_9595_), .C(_9321_), .Y(_9625_) );
	OAI21X1 OAI21X1_4046 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9624_), .C(_9625_), .Y(_9626_) );
	OAI21X1 OAI21X1_4047 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9285__bF_buf2), .C(_9149__bF_buf3), .Y(_9627_) );
	AOI21X1 AOI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_13_), .B(_9326_), .C(_9627_), .Y(_9628_) );
	NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_9628_), .B(_9626_), .Y(_9629_) );
	AOI22X1 AOI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(_8861__bF_buf0), .B(_9629_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf3), .D(_9621_), .Y(_9630_) );
	OAI21X1 OAI21X1_4048 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .B(_9149__bF_buf2), .C(_9251__bF_buf3), .Y(_9631_) );
	AOI21X1 AOI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(csr_gpr_iu_csr_pc_next_12_), .C(_9094__bF_buf5), .Y(_9632_) );
	OAI21X1 OAI21X1_4049 ( .gnd(gnd), .vdd(vdd), .A(_9631_), .B(_9630_), .C(_9632_), .Y(_9633_) );
	OAI22X1 OAI22X1_755 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(biu_mmu_msu_0_bF_buf4), .C(_8912_), .D(_9105__bF_buf0), .Y(_9634_) );
	AOI21X1 AOI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_12_), .B(_9098__bF_buf0), .C(_9634_), .Y(_9635_) );
	AOI21X1 AOI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_9635_), .B(_9094__bF_buf4), .C(_7303__bF_buf10_bF_buf0), .Y(_9636_) );
	NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_9636_), .B(_9633_), .Y(_9637_) );
	AOI21X1 AOI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_9637_), .B(_9614_), .C(rst_bF_buf35), .Y(_6725__12_) );
	INVX1 INVX1_1641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_13_), .Y(_9638_) );
	AOI21X1 AOI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf0), .B(_9638_), .C(_7304__bF_buf6_bF_buf0), .Y(_9639_) );
	OAI21X1 OAI21X1_4050 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(_9268__bF_buf6), .C(_9639_), .Y(_9640_) );
	NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_11_), .B(_9575_), .Y(_9641_) );
	OAI21X1 OAI21X1_4051 ( .gnd(gnd), .vdd(vdd), .A(_9615_), .B(_9641_), .C(_9049_), .Y(_9642_) );
	NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_9615_), .B(_9049_), .Y(_9643_) );
	INVX1 INVX1_1642 ( .gnd(gnd), .vdd(vdd), .A(_9643_), .Y(_9644_) );
	OAI21X1 OAI21X1_4052 ( .gnd(gnd), .vdd(vdd), .A(_9641_), .B(_9644_), .C(_9642_), .Y(_9645_) );
	AOI22X1 AOI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_13_), .B(_9273__bF_buf1), .C(csr_gpr_iu_csr_mtvec_14_), .D(_9281__bF_buf0), .Y(_9646_) );
	OAI21X1 OAI21X1_4053 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_9645_), .C(_9646_), .Y(_9647_) );
	NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_9647_), .Y(_9648_) );
	OAI21X1 OAI21X1_4054 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7742_), .C(_7427_), .Y(_9649_) );
	NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9624_), .Y(_9650_) );
	NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_13_), .B(_9650_), .Y(_9651_) );
	NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_12_), .B(csr_gpr_iu_csr_stvec_13_), .Y(_9652_) );
	OAI21X1 OAI21X1_4055 ( .gnd(gnd), .vdd(vdd), .A(_9652_), .B(_9624_), .C(_9322__bF_buf2), .Y(_9653_) );
	OAI21X1 OAI21X1_4056 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .B(_9285__bF_buf1), .C(_7426_), .Y(_9654_) );
	AOI21X1 AOI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_14_), .B(_9326_), .C(_9654_), .Y(_9655_) );
	OAI21X1 OAI21X1_4057 ( .gnd(gnd), .vdd(vdd), .A(_9653_), .B(_9651_), .C(_9655_), .Y(_9656_) );
	AOI21X1 AOI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_9656_), .B(_9649_), .C(_7424__bF_buf1), .Y(_9657_) );
	OAI21X1 OAI21X1_4058 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(_7423_), .C(_9251__bF_buf2), .Y(_9658_) );
	AOI21X1 AOI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_9648_), .B(_9657_), .C(_9658_), .Y(_9659_) );
	OAI21X1 OAI21X1_4059 ( .gnd(gnd), .vdd(vdd), .A(_9638_), .B(_9251__bF_buf1), .C(_9095__bF_buf4), .Y(_9660_) );
	OAI22X1 OAI22X1_756 ( .gnd(gnd), .vdd(vdd), .A(_7742_), .B(biu_mmu_msu_0_bF_buf3), .C(_8918_), .D(_9105__bF_buf4), .Y(_9661_) );
	AOI21X1 AOI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_13_), .B(_9098__bF_buf4), .C(_9661_), .Y(_9662_) );
	AOI21X1 AOI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_9662_), .B(_9094__bF_buf3), .C(_7303__bF_buf9_bF_buf0), .Y(_9663_) );
	OAI21X1 OAI21X1_4060 ( .gnd(gnd), .vdd(vdd), .A(_9660_), .B(_9659_), .C(_9663_), .Y(_9664_) );
	AOI21X1 AOI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_9664_), .B(_9640_), .C(rst_bF_buf34), .Y(_6725__13_) );
	INVX1 INVX1_1643 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_14_), .Y(_9665_) );
	AOI21X1 AOI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf5), .B(_9665_), .C(_7304__bF_buf5), .Y(_9666_) );
	OAI21X1 OAI21X1_4061 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(_9268__bF_buf4), .C(_9666_), .Y(_9667_) );
	OAI21X1 OAI21X1_4062 ( .gnd(gnd), .vdd(vdd), .A(_9644_), .B(_9641_), .C(csr_gpr_iu_csr_mtvec_14_), .Y(_9668_) );
	INVX1 INVX1_1644 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_14_), .Y(_9669_) );
	NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_9669_), .B(_9643_), .C(_9617_), .Y(_9670_) );
	AOI21X1 AOI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_9670_), .B(_9668_), .C(_9275_), .Y(_9671_) );
	OAI22X1 OAI22X1_757 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_9280_), .C(_9669_), .D(_9274_), .Y(_9672_) );
	OAI21X1 OAI21X1_4063 ( .gnd(gnd), .vdd(vdd), .A(_9672_), .B(_9671_), .C(_8614_), .Y(_9673_) );
	OAI21X1 OAI21X1_4064 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7755_), .C(_7427_), .Y(_9674_) );
	NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_9652_), .B(_9624_), .Y(_9675_) );
	AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_9675_), .B(csr_gpr_iu_csr_stvec_14_), .Y(_9676_) );
	OAI21X1 OAI21X1_4065 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_14_), .B(_9675_), .C(_9322__bF_buf1), .Y(_9677_) );
	INVX1 INVX1_1645 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_14_), .Y(_9678_) );
	OAI21X1 OAI21X1_4066 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_9285__bF_buf0), .C(_7426_), .Y(_9679_) );
	AOI21X1 AOI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_15_), .B(_9326_), .C(_9679_), .Y(_9680_) );
	OAI21X1 OAI21X1_4067 ( .gnd(gnd), .vdd(vdd), .A(_9676_), .B(_9677_), .C(_9680_), .Y(_9681_) );
	AOI21X1 AOI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_9681_), .B(_9674_), .C(_7424__bF_buf0), .Y(_9682_) );
	OAI21X1 OAI21X1_4068 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(_7423_), .C(_9251__bF_buf0), .Y(_9683_) );
	AOI21X1 AOI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_9673_), .B(_9682_), .C(_9683_), .Y(_9684_) );
	OAI21X1 OAI21X1_4069 ( .gnd(gnd), .vdd(vdd), .A(_9665_), .B(_9251__bF_buf6), .C(_9095__bF_buf3), .Y(_9685_) );
	OAI22X1 OAI22X1_758 ( .gnd(gnd), .vdd(vdd), .A(_7755_), .B(biu_mmu_msu_0_bF_buf2), .C(_8927_), .D(_9105__bF_buf3), .Y(_9686_) );
	AOI21X1 AOI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_14_), .B(_9098__bF_buf3), .C(_9686_), .Y(_9687_) );
	AOI21X1 AOI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_9687_), .B(_9094__bF_buf2), .C(_7303__bF_buf8_bF_buf0), .Y(_9688_) );
	OAI21X1 OAI21X1_4070 ( .gnd(gnd), .vdd(vdd), .A(_9685_), .B(_9684_), .C(_9688_), .Y(_9689_) );
	AOI21X1 AOI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_9689_), .B(_9667_), .C(rst_bF_buf33), .Y(_6725__14_) );
	INVX1 INVX1_1646 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_15_), .Y(_9690_) );
	AOI21X1 AOI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf3), .B(_9690_), .C(_7304__bF_buf4), .Y(_9691_) );
	OAI21X1 OAI21X1_4071 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .B(_9268__bF_buf2), .C(_9691_), .Y(_9692_) );
	NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_14_), .B(_9643_), .C(_9617_), .Y(_9693_) );
	NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_9545_), .B(_9600_), .Y(_9694_) );
	AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_9572_), .B(_9694_), .Y(_9695_) );
	NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_14_), .B(csr_gpr_iu_csr_mtvec_15_), .Y(_9696_) );
	NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_9696_), .B(_9644_), .Y(_9697_) );
	NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_9694_), .B(_9571_), .C(_9697_), .Y(_9698_) );
	INVX1 INVX1_1647 ( .gnd(gnd), .vdd(vdd), .A(_9698_), .Y(_9699_) );
	AOI22X1 AOI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(_9695_), .B(_9697_), .C(_9699_), .D(_9503_), .Y(_9700_) );
	NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf0), .B(_9700_), .Y(_9701_) );
	AOI21X1 AOI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_9693_), .B(_9053_), .C(_9701_), .Y(_9702_) );
	INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_16_), .Y(_9703_) );
	OAI22X1 OAI22X1_759 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9280_), .C(_9053_), .D(_9274_), .Y(_9704_) );
	OAI21X1 OAI21X1_4072 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9702_), .C(_8614_), .Y(_9705_) );
	OAI21X1 OAI21X1_4073 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7766_), .C(_7427_), .Y(_9706_) );
	AOI21X1 AOI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_9675_), .B(csr_gpr_iu_csr_stvec_14_), .C(csr_gpr_iu_csr_stvec_15_), .Y(_9707_) );
	AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .B(_9623_), .Y(_9708_) );
	NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_14_), .B(csr_gpr_iu_csr_stvec_15_), .Y(_9709_) );
	NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_9652_), .B(_9709_), .Y(_9710_) );
	NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9710_), .C(_9560_), .Y(_9711_) );
	INVX1 INVX1_1648 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .Y(_9712_) );
	AOI22X1 AOI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(_9708_), .B(_9710_), .C(_9712_), .D(_9488_), .Y(_9713_) );
	NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf0), .B(_9713_), .Y(_9714_) );
	OAI21X1 OAI21X1_4074 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_9285__bF_buf4), .C(_7426_), .Y(_9715_) );
	AOI21X1 AOI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_16_), .B(_9326_), .C(_9715_), .Y(_9716_) );
	OAI21X1 OAI21X1_4075 ( .gnd(gnd), .vdd(vdd), .A(_9714_), .B(_9707_), .C(_9716_), .Y(_9717_) );
	AOI21X1 AOI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_9717_), .B(_9706_), .C(_7424__bF_buf3), .Y(_9718_) );
	OAI21X1 OAI21X1_4076 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .B(_7423_), .C(_9251__bF_buf5), .Y(_9719_) );
	AOI21X1 AOI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .B(_9718_), .C(_9719_), .Y(_9720_) );
	OAI21X1 OAI21X1_4077 ( .gnd(gnd), .vdd(vdd), .A(_9690_), .B(_9251__bF_buf4), .C(_9095__bF_buf2), .Y(_9721_) );
	OAI22X1 OAI22X1_760 ( .gnd(gnd), .vdd(vdd), .A(_7766_), .B(biu_mmu_msu_0_bF_buf1), .C(_8930_), .D(_9105__bF_buf2), .Y(_9722_) );
	AOI21X1 AOI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_15_), .B(_9098__bF_buf2), .C(_9722_), .Y(_9723_) );
	AOI21X1 AOI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_9723_), .B(_9094__bF_buf1), .C(_7303__bF_buf7_bF_buf0), .Y(_9724_) );
	OAI21X1 OAI21X1_4078 ( .gnd(gnd), .vdd(vdd), .A(_9721_), .B(_9720_), .C(_9724_), .Y(_9725_) );
	AOI21X1 AOI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_9725_), .B(_9692_), .C(rst_bF_buf32), .Y(_6725__15_) );
	INVX1 INVX1_1649 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .Y(_9726_) );
	OAI21X1 OAI21X1_4079 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9246_), .C(csr_gpr_iu_csr_pc_next_16_), .Y(_9727_) );
	OAI21X1 OAI21X1_4080 ( .gnd(gnd), .vdd(vdd), .A(_9726_), .B(_9268__bF_buf1), .C(_9727_), .Y(_9728_) );
	NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6_bF_buf0), .B(_9728_), .Y(_9729_) );
	INVX1 INVX1_1650 ( .gnd(gnd), .vdd(vdd), .A(_9700_), .Y(_9730_) );
	NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_16_), .B(_9730_), .Y(_9731_) );
	OAI21X1 OAI21X1_4081 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9700_), .C(_9276__bF_buf3), .Y(_9732_) );
	AOI22X1 AOI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_16_), .B(_9273__bF_buf0), .C(csr_gpr_iu_csr_mtvec_17_), .D(_9281__bF_buf3), .Y(_9733_) );
	OAI21X1 OAI21X1_4082 ( .gnd(gnd), .vdd(vdd), .A(_9732_), .B(_9731_), .C(_9733_), .Y(_9734_) );
	INVX1 INVX1_1651 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_16_), .Y(_9735_) );
	AOI21X1 AOI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_9713_), .B(_9735_), .C(_9321_), .Y(_9736_) );
	OAI21X1 OAI21X1_4083 ( .gnd(gnd), .vdd(vdd), .A(_9735_), .B(_9713_), .C(_9736_), .Y(_9737_) );
	OAI21X1 OAI21X1_4084 ( .gnd(gnd), .vdd(vdd), .A(_9735_), .B(_9285__bF_buf3), .C(_9149__bF_buf1), .Y(_9738_) );
	AOI21X1 AOI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_17_), .B(_9326_), .C(_9738_), .Y(_9739_) );
	NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_9739_), .B(_9737_), .Y(_9740_) );
	AOI22X1 AOI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf2), .B(_9734_), .C(_8861__bF_buf6), .D(_9740_), .Y(_9741_) );
	OAI21X1 OAI21X1_4085 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .B(_9149__bF_buf0), .C(_9251__bF_buf3), .Y(_9742_) );
	AOI21X1 AOI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(csr_gpr_iu_csr_pc_next_16_), .C(_9094__bF_buf0), .Y(_9743_) );
	OAI21X1 OAI21X1_4086 ( .gnd(gnd), .vdd(vdd), .A(_9742_), .B(_9741_), .C(_9743_), .Y(_9744_) );
	OAI22X1 OAI22X1_761 ( .gnd(gnd), .vdd(vdd), .A(_9726_), .B(biu_mmu_msu_0_bF_buf0), .C(_8935_), .D(_9105__bF_buf1), .Y(_9745_) );
	AOI21X1 AOI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_16_), .B(_9098__bF_buf1), .C(_9745_), .Y(_9746_) );
	AOI21X1 AOI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_9746_), .B(_9094__bF_buf5), .C(_7303__bF_buf5_bF_buf0), .Y(_9747_) );
	NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_9747_), .B(_9744_), .Y(_9748_) );
	AOI21X1 AOI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_9729_), .B(_9748_), .C(rst_bF_buf31), .Y(_6725__16_) );
	INVX1 INVX1_1652 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_17_), .Y(_9749_) );
	AOI21X1 AOI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf0), .B(_9749_), .C(_7304__bF_buf3), .Y(_9750_) );
	OAI21X1 OAI21X1_4087 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(_9268__bF_buf6), .C(_9750_), .Y(_9751_) );
	OAI21X1 OAI21X1_4088 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9700_), .C(_9057_), .Y(_9752_) );
	NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_16_), .B(csr_gpr_iu_csr_mtvec_17_), .Y(_9753_) );
	OAI21X1 OAI21X1_4089 ( .gnd(gnd), .vdd(vdd), .A(_9700_), .B(_9753_), .C(_9752_), .Y(_9754_) );
	OAI21X1 OAI21X1_4090 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_9274_), .C(_8614_), .Y(_9755_) );
	AOI21X1 AOI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(_9281__bF_buf2), .C(_9755_), .Y(_9756_) );
	OAI21X1 OAI21X1_4091 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_9754_), .C(_9756_), .Y(_9757_) );
	NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9710_), .C(_9562_), .Y(_9758_) );
	OAI21X1 OAI21X1_4092 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .B(_9527_), .C(_9758_), .Y(_9759_) );
	AOI21X1 AOI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_9759_), .B(csr_gpr_iu_csr_stvec_16_), .C(csr_gpr_iu_csr_stvec_17_), .Y(_9760_) );
	NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_16_), .B(csr_gpr_iu_csr_stvec_17_), .Y(_9761_) );
	OAI21X1 OAI21X1_4093 ( .gnd(gnd), .vdd(vdd), .A(_9761_), .B(_9713_), .C(_9322__bF_buf3), .Y(_9762_) );
	OAI21X1 OAI21X1_4094 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_9285__bF_buf2), .C(_7426_), .Y(_9763_) );
	AOI21X1 AOI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_18_), .B(_9326_), .C(_9763_), .Y(_9764_) );
	OAI21X1 OAI21X1_4095 ( .gnd(gnd), .vdd(vdd), .A(_9762_), .B(_9760_), .C(_9764_), .Y(_9765_) );
	AOI21X1 AOI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7787_), .C(_7424__bF_buf2), .Y(_9766_) );
	NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_9766_), .B(_9765_), .C(_9757_), .Y(_9767_) );
	OAI21X1 OAI21X1_4096 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .B(_7423_), .C(_9767_), .Y(_9768_) );
	NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_9251__bF_buf2), .B(_9768_), .Y(_9769_) );
	OAI21X1 OAI21X1_4097 ( .gnd(gnd), .vdd(vdd), .A(_9749_), .B(_9251__bF_buf1), .C(_9769_), .Y(_9770_) );
	OAI22X1 OAI22X1_762 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .B(biu_mmu_msu_0_bF_buf4), .C(_8941_), .D(_9105__bF_buf0), .Y(_9771_) );
	AOI21X1 AOI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_17_), .B(_9098__bF_buf0), .C(_9771_), .Y(_9772_) );
	AOI21X1 AOI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_9772_), .B(_9094__bF_buf4), .C(_7303__bF_buf4_bF_buf0), .Y(_9773_) );
	OAI21X1 OAI21X1_4098 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf3), .B(_9770_), .C(_9773_), .Y(_9774_) );
	AOI21X1 AOI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_9774_), .B(_9751_), .C(rst_bF_buf30), .Y(_6725__17_) );
	INVX1 INVX1_1653 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_18_), .Y(_9775_) );
	AOI21X1 AOI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf5), .B(_9775_), .C(_7304__bF_buf2), .Y(_9776_) );
	OAI21X1 OAI21X1_4099 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(_9268__bF_buf4), .C(_9776_), .Y(_9777_) );
	NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_9753_), .B(_9700_), .Y(_9778_) );
	NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(_9778_), .Y(_9779_) );
	NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(_9778_), .Y(_9780_) );
	NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf2), .B(_9780_), .Y(_9781_) );
	AOI22X1 AOI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(_9273__bF_buf3), .C(csr_gpr_iu_csr_mtvec_19_), .D(_9281__bF_buf1), .Y(_9782_) );
	OAI21X1 OAI21X1_4100 ( .gnd(gnd), .vdd(vdd), .A(_9779_), .B(_9781_), .C(_9782_), .Y(_9783_) );
	NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf1), .B(_9783_), .Y(_9784_) );
	INVX1 INVX1_1654 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_18_), .Y(_9785_) );
	NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_16_), .B(csr_gpr_iu_csr_stvec_17_), .C(_9759_), .Y(_9786_) );
	OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_9786_), .B(_9785_), .Y(_9787_) );
	AOI21X1 AOI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_9786_), .B(_9785_), .C(_9321_), .Y(_9788_) );
	AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_9787_), .B(_9788_), .Y(_9789_) );
	AOI21X1 AOI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_18_), .B(_9284_), .C(_9291_), .Y(_9790_) );
	OAI21X1 OAI21X1_4101 ( .gnd(gnd), .vdd(vdd), .A(_8086_), .B(_9325_), .C(_9790_), .Y(_9791_) );
	OAI21X1 OAI21X1_4102 ( .gnd(gnd), .vdd(vdd), .A(_9791_), .B(_9789_), .C(_8861__bF_buf5), .Y(_9792_) );
	OAI21X1 OAI21X1_4103 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(_9149__bF_buf4), .C(_9251__bF_buf0), .Y(_9793_) );
	AOI21X1 AOI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_9784_), .B(_9792_), .C(_9793_), .Y(_9794_) );
	OAI21X1 OAI21X1_4104 ( .gnd(gnd), .vdd(vdd), .A(_9775_), .B(_9251__bF_buf6), .C(_9095__bF_buf1), .Y(_9795_) );
	OAI22X1 OAI22X1_763 ( .gnd(gnd), .vdd(vdd), .A(_7800_), .B(biu_mmu_msu_0_bF_buf3), .C(_8947_), .D(_9105__bF_buf4), .Y(_9796_) );
	AOI21X1 AOI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_18_), .B(_9098__bF_buf4), .C(_9796_), .Y(_9797_) );
	AOI21X1 AOI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_9797_), .B(_9094__bF_buf2), .C(_7303__bF_buf3_bF_buf0), .Y(_9798_) );
	OAI21X1 OAI21X1_4105 ( .gnd(gnd), .vdd(vdd), .A(_9795_), .B(_9794_), .C(_9798_), .Y(_9799_) );
	AOI21X1 AOI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_9799_), .B(_9777_), .C(rst_bF_buf29), .Y(_6725__18_) );
	INVX1 INVX1_1655 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_19_), .Y(_9800_) );
	AOI21X1 AOI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf3), .B(_9800_), .C(_7304__bF_buf1), .Y(_9801_) );
	OAI21X1 OAI21X1_4106 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .B(_9268__bF_buf2), .C(_9801_), .Y(_9802_) );
	NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_18_), .B(csr_gpr_iu_csr_stvec_19_), .Y(_9803_) );
	NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_9761_), .B(_9803_), .Y(_9804_) );
	INVX1 INVX1_1656 ( .gnd(gnd), .vdd(vdd), .A(_9804_), .Y(_9805_) );
	OAI21X1 OAI21X1_4107 ( .gnd(gnd), .vdd(vdd), .A(_9805_), .B(_9713_), .C(_9322__bF_buf2), .Y(_9806_) );
	AOI21X1 AOI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_9787_), .B(_8086_), .C(_9806_), .Y(_9807_) );
	INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_20_), .Y(_9808_) );
	AOI21X1 AOI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_19_), .B(_9284_), .C(_9291_), .Y(_9809_) );
	OAI21X1 OAI21X1_4108 ( .gnd(gnd), .vdd(vdd), .A(_9808_), .B(_9325_), .C(_9809_), .Y(_9810_) );
	OAI21X1 OAI21X1_4109 ( .gnd(gnd), .vdd(vdd), .A(_9810_), .B(_9807_), .C(_8861__bF_buf4), .Y(_9811_) );
	NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_9274_), .Y(_9812_) );
	OAI21X1 OAI21X1_4110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_31_), .B(csr_gpr_iu_csr_mtvec_20_), .C(_9274_), .Y(_9813_) );
	NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_9780_), .Y(_9814_) );
	NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(csr_gpr_iu_csr_mtvec_19_), .C(_9778_), .Y(_9815_) );
	NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_9815_), .B(_9814_), .Y(_9816_) );
	AOI21X1 AOI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_9816_), .B(csr_gpr_iu_csr_mcause_31_), .C(_9813_), .Y(_9817_) );
	OAI21X1 OAI21X1_4111 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .B(_9817_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf0), .Y(_9818_) );
	OAI21X1 OAI21X1_4112 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .B(_9149__bF_buf3), .C(_9251__bF_buf5), .Y(_9819_) );
	AOI21X1 AOI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_9818_), .B(_9811_), .C(_9819_), .Y(_9820_) );
	OAI21X1 OAI21X1_4113 ( .gnd(gnd), .vdd(vdd), .A(_9800_), .B(_9251__bF_buf4), .C(_9095__bF_buf0), .Y(_9821_) );
	OAI22X1 OAI22X1_764 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .B(biu_mmu_msu_0_bF_buf2), .C(_8952_), .D(_9105__bF_buf3), .Y(_9822_) );
	AOI21X1 AOI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_19_), .B(_9098__bF_buf3), .C(_9822_), .Y(_9823_) );
	AOI21X1 AOI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_9823_), .B(_9094__bF_buf1), .C(_7303__bF_buf2), .Y(_9824_) );
	OAI21X1 OAI21X1_4114 ( .gnd(gnd), .vdd(vdd), .A(_9821_), .B(_9820_), .C(_9824_), .Y(_9825_) );
	AOI21X1 AOI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .B(_9802_), .C(rst_bF_buf28), .Y(_6725__19_) );
	INVX1 INVX1_1657 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_20_), .Y(_9826_) );
	AOI21X1 AOI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf1), .B(_9826_), .C(_7304__bF_buf0), .Y(_9827_) );
	OAI21X1 OAI21X1_4115 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_9268__bF_buf0), .C(_9827_), .Y(_9828_) );
	NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(csr_gpr_iu_csr_mtvec_19_), .Y(_9829_) );
	NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_9753_), .B(_9829_), .Y(_9830_) );
	INVX1 INVX1_1658 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .Y(_9831_) );
	NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_9831_), .B(_9700_), .Y(_9832_) );
	NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_20_), .B(_9832_), .Y(_9833_) );
	NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_20_), .B(_9832_), .Y(_9834_) );
	NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf1), .B(_9834_), .Y(_9835_) );
	AOI22X1 AOI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_20_), .B(_9273__bF_buf2), .C(csr_gpr_iu_csr_mtvec_21_), .D(_9281__bF_buf0), .Y(_9836_) );
	OAI21X1 OAI21X1_4116 ( .gnd(gnd), .vdd(vdd), .A(_9833_), .B(_9835_), .C(_9836_), .Y(_9837_) );
	NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_1_bF_buf3), .B(_9837_), .Y(_9838_) );
	OAI21X1 OAI21X1_4117 ( .gnd(gnd), .vdd(vdd), .A(_9808_), .B(_9285__bF_buf1), .C(_9149__bF_buf2), .Y(_9839_) );
	AOI21X1 AOI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_9487_), .C(_9711_), .Y(_9840_) );
	INVX1 INVX1_1659 ( .gnd(gnd), .vdd(vdd), .A(_9758_), .Y(_9841_) );
	OAI21X1 OAI21X1_4118 ( .gnd(gnd), .vdd(vdd), .A(_9841_), .B(_9840_), .C(_9804_), .Y(_9842_) );
	OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_9842_), .B(_9808_), .Y(_9843_) );
	OAI21X1 OAI21X1_4119 ( .gnd(gnd), .vdd(vdd), .A(_9805_), .B(_9713_), .C(_9808_), .Y(_9844_) );
	NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_9844_), .B(_9843_), .Y(_9845_) );
	OAI21X1 OAI21X1_4120 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf0), .B(csr_gpr_iu_csr_stvec_21_), .C(_9285__bF_buf0), .Y(_9846_) );
	AOI21X1 AOI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_9845_), .B(csr_gpr_iu_csr_scause_31_bF_buf3), .C(_9846_), .Y(_9847_) );
	OAI21X1 OAI21X1_4121 ( .gnd(gnd), .vdd(vdd), .A(_9839_), .B(_9847_), .C(_8861__bF_buf3), .Y(_9848_) );
	OAI21X1 OAI21X1_4122 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_9149__bF_buf1), .C(_9251__bF_buf3), .Y(_9849_) );
	AOI21X1 AOI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_9848_), .B(_9838_), .C(_9849_), .Y(_9850_) );
	OAI21X1 OAI21X1_4123 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .B(_9251__bF_buf2), .C(_9095__bF_buf4), .Y(_9851_) );
	NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_9097_), .Y(_9852_) );
	OAI21X1 OAI21X1_4124 ( .gnd(gnd), .vdd(vdd), .A(_8957_), .B(_9105__bF_buf2), .C(_9852_), .Y(_9853_) );
	AOI21X1 AOI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_20_), .B(_9098__bF_buf2), .C(_9853_), .Y(_9854_) );
	AOI21X1 AOI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_9854_), .B(_9094__bF_buf0), .C(_7303__bF_buf1), .Y(_9855_) );
	OAI21X1 OAI21X1_4125 ( .gnd(gnd), .vdd(vdd), .A(_9851_), .B(_9850_), .C(_9855_), .Y(_9856_) );
	AOI21X1 AOI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_9856_), .B(_9828_), .C(rst_bF_buf27), .Y(_6725__20_) );
	INVX1 INVX1_1660 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_21_), .Y(_9857_) );
	AOI21X1 AOI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf6), .B(_9857_), .C(_7304__bF_buf14_bF_buf3), .Y(_9858_) );
	OAI21X1 OAI21X1_4126 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .B(_9268__bF_buf5), .C(_9858_), .Y(_9859_) );
	AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_9832_), .B(csr_gpr_iu_csr_mtvec_20_), .Y(_9860_) );
	NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_21_), .B(_9860_), .Y(_9861_) );
	OAI21X1 OAI21X1_4127 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9834_), .C(_9276__bF_buf0), .Y(_9862_) );
	OAI21X1 OAI21X1_4128 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9274_), .C(_8614_), .Y(_9863_) );
	AOI21X1 AOI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_22_), .B(_9281__bF_buf3), .C(_9863_), .Y(_9864_) );
	OAI21X1 OAI21X1_4129 ( .gnd(gnd), .vdd(vdd), .A(_9862_), .B(_9861_), .C(_9864_), .Y(_9865_) );
	AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .B(_8089_), .Y(_9866_) );
	OAI21X1 OAI21X1_4130 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .B(_9843_), .C(_9322__bF_buf1), .Y(_9867_) );
	OAI21X1 OAI21X1_4131 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .B(_9285__bF_buf4), .C(_7426_), .Y(_9868_) );
	AOI21X1 AOI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_22_), .B(_9326_), .C(_9868_), .Y(_9869_) );
	OAI21X1 OAI21X1_4132 ( .gnd(gnd), .vdd(vdd), .A(_9866_), .B(_9867_), .C(_9869_), .Y(_9870_) );
	AOI21X1 AOI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7840_), .C(_7424__bF_buf1), .Y(_9871_) );
	NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_9870_), .B(_9871_), .C(_9865_), .Y(_9872_) );
	AOI21X1 AOI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .B(_7424__bF_buf0), .C(_9292_), .Y(_9873_) );
	AOI22X1 AOI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(_9857_), .B(_9292_), .C(_9873_), .D(_9872_), .Y(_9874_) );
	OAI22X1 OAI22X1_765 ( .gnd(gnd), .vdd(vdd), .A(_7840_), .B(biu_mmu_msu_0_bF_buf1), .C(_8962_), .D(_9105__bF_buf1), .Y(_9875_) );
	AOI21X1 AOI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_21_), .B(_9098__bF_buf1), .C(_9875_), .Y(_9876_) );
	AOI21X1 AOI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_9876_), .B(_9094__bF_buf5), .C(_7303__bF_buf0), .Y(_9877_) );
	OAI21X1 OAI21X1_4133 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf4), .B(_9874_), .C(_9877_), .Y(_9878_) );
	AOI21X1 AOI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_9878_), .B(_9859_), .C(rst_bF_buf26), .Y(_6725__21_) );
	INVX1 INVX1_1661 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_22_), .Y(_9879_) );
	AOI21X1 AOI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf4), .B(_9879_), .C(_7304__bF_buf13_bF_buf3), .Y(_9880_) );
	OAI21X1 OAI21X1_4134 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_9268__bF_buf3), .C(_9880_), .Y(_9881_) );
	OAI21X1 OAI21X1_4135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7839_), .C(_7427_), .Y(_9882_) );
	INVX1 INVX1_1662 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .Y(_9883_) );
	AOI21X1 AOI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_9883_), .B(csr_gpr_iu_csr_stvec_21_), .C(csr_gpr_iu_csr_stvec_22_), .Y(_9884_) );
	NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_21_), .B(csr_gpr_iu_csr_stvec_22_), .Y(_9885_) );
	OAI21X1 OAI21X1_4136 ( .gnd(gnd), .vdd(vdd), .A(_9885_), .B(_9843_), .C(_9322__bF_buf0), .Y(_9886_) );
	NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_9886_), .B(_9884_), .Y(_9887_) );
	AOI21X1 AOI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_22_), .B(_9284_), .C(_7427_), .Y(_9888_) );
	OAI21X1 OAI21X1_4137 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_9325_), .C(_9888_), .Y(_9889_) );
	OAI21X1 OAI21X1_4138 ( .gnd(gnd), .vdd(vdd), .A(_9889_), .B(_9887_), .C(_9882_), .Y(_9890_) );
	AOI21X1 AOI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_9860_), .B(csr_gpr_iu_csr_mtvec_21_), .C(csr_gpr_iu_csr_mtvec_22_), .Y(_9891_) );
	NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_21_), .B(csr_gpr_iu_csr_mtvec_22_), .Y(_9892_) );
	OAI21X1 OAI21X1_4139 ( .gnd(gnd), .vdd(vdd), .A(_9892_), .B(_9834_), .C(_9276__bF_buf3), .Y(_9893_) );
	AOI22X1 AOI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_22_), .B(_9273__bF_buf1), .C(csr_gpr_iu_csr_mtvec_23_), .D(_9281__bF_buf2), .Y(_9894_) );
	OAI21X1 OAI21X1_4140 ( .gnd(gnd), .vdd(vdd), .A(_9893_), .B(_9891_), .C(_9894_), .Y(_9895_) );
	AOI21X1 AOI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_9895_), .B(_8614_), .C(_7424__bF_buf3), .Y(_9896_) );
	OAI21X1 OAI21X1_4141 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_7423_), .C(_9251__bF_buf1), .Y(_9897_) );
	AOI21X1 AOI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_9896_), .B(_9890_), .C(_9897_), .Y(_9898_) );
	OAI21X1 OAI21X1_4142 ( .gnd(gnd), .vdd(vdd), .A(_9879_), .B(_9251__bF_buf0), .C(_9095__bF_buf3), .Y(_9899_) );
	OAI22X1 OAI22X1_766 ( .gnd(gnd), .vdd(vdd), .A(_7839_), .B(biu_mmu_msu_0_bF_buf0), .C(_8967_), .D(_9105__bF_buf0), .Y(_9900_) );
	AOI21X1 AOI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_22_), .B(_9098__bF_buf0), .C(_9900_), .Y(_9901_) );
	AOI21X1 AOI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_9901_), .B(_9094__bF_buf3), .C(_7303__bF_buf14_bF_buf3), .Y(_9902_) );
	OAI21X1 OAI21X1_4143 ( .gnd(gnd), .vdd(vdd), .A(_9899_), .B(_9898_), .C(_9902_), .Y(_9903_) );
	AOI21X1 AOI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_9903_), .B(_9881_), .C(rst_bF_buf25), .Y(_6725__22_) );
	INVX1 INVX1_1663 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_23_), .Y(_9904_) );
	AOI21X1 AOI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf2), .B(_9904_), .C(_7304__bF_buf12_bF_buf3), .Y(_9905_) );
	OAI21X1 OAI21X1_4144 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .B(_9268__bF_buf1), .C(_9905_), .Y(_9906_) );
	OAI21X1 OAI21X1_4145 ( .gnd(gnd), .vdd(vdd), .A(_9885_), .B(_9843_), .C(_8092_), .Y(_9907_) );
	NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_20_), .B(csr_gpr_iu_csr_stvec_21_), .Y(_9908_) );
	NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_22_), .B(csr_gpr_iu_csr_stvec_23_), .Y(_9909_) );
	NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_9908_), .B(_9909_), .Y(_9910_) );
	NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_9804_), .B(_9910_), .Y(_9911_) );
	INVX1 INVX1_1664 ( .gnd(gnd), .vdd(vdd), .A(_9911_), .Y(_9912_) );
	OAI21X1 OAI21X1_4146 ( .gnd(gnd), .vdd(vdd), .A(_9841_), .B(_9840_), .C(_9912_), .Y(_9913_) );
	INVX1 INVX1_1665 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9914_) );
	NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_9914_), .Y(_9915_) );
	AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_9907_), .B(_9915_), .Y(_9916_) );
	INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_24_), .Y(_9917_) );
	AOI21X1 AOI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_23_), .B(_9284_), .C(_9291_), .Y(_9918_) );
	OAI21X1 OAI21X1_4147 ( .gnd(gnd), .vdd(vdd), .A(_9917_), .B(_9325_), .C(_9918_), .Y(_9919_) );
	OAI21X1 OAI21X1_4148 ( .gnd(gnd), .vdd(vdd), .A(_9919_), .B(_9916_), .C(_8861__bF_buf2), .Y(_9920_) );
	OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_9834_), .B(_9892_), .Y(_9921_) );
	OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_9892_), .B(_9069_), .Y(_9922_) );
	OAI21X1 OAI21X1_4149 ( .gnd(gnd), .vdd(vdd), .A(_9922_), .B(_9834_), .C(_9276__bF_buf2), .Y(_9923_) );
	AOI21X1 AOI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_9921_), .B(_9069_), .C(_9923_), .Y(_9924_) );
	INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_24_), .Y(_9925_) );
	OAI22X1 OAI22X1_767 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9280_), .C(_9069_), .D(_9274_), .Y(_9926_) );
	OAI21X1 OAI21X1_4150 ( .gnd(gnd), .vdd(vdd), .A(_9926_), .B(_9924_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf2), .Y(_9927_) );
	OAI21X1 OAI21X1_4151 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .B(_9149__bF_buf0), .C(_9251__bF_buf6), .Y(_9928_) );
	AOI21X1 AOI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_9927_), .B(_9920_), .C(_9928_), .Y(_9929_) );
	OAI21X1 OAI21X1_4152 ( .gnd(gnd), .vdd(vdd), .A(_9904_), .B(_9251__bF_buf5), .C(_9095__bF_buf2), .Y(_9930_) );
	OAI22X1 OAI22X1_768 ( .gnd(gnd), .vdd(vdd), .A(_7850_), .B(biu_mmu_msu_0_bF_buf4), .C(_8972_), .D(_9105__bF_buf4), .Y(_9931_) );
	AOI21X1 AOI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_23_), .B(_9098__bF_buf4), .C(_9931_), .Y(_9932_) );
	AOI21X1 AOI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_9094__bF_buf2), .C(_7303__bF_buf13_bF_buf3), .Y(_9933_) );
	OAI21X1 OAI21X1_4153 ( .gnd(gnd), .vdd(vdd), .A(_9930_), .B(_9929_), .C(_9933_), .Y(_9934_) );
	AOI21X1 AOI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_9906_), .C(rst_bF_buf24), .Y(_6725__23_) );
	INVX1 INVX1_1666 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_24_), .Y(_9935_) );
	AOI21X1 AOI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf0), .B(_9935_), .C(_7304__bF_buf11_bF_buf3), .Y(_9936_) );
	OAI21X1 OAI21X1_4154 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .B(_9268__bF_buf6), .C(_9936_), .Y(_9937_) );
	NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_20_), .B(csr_gpr_iu_csr_mtvec_21_), .Y(_9938_) );
	NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_22_), .B(csr_gpr_iu_csr_mtvec_23_), .Y(_9939_) );
	NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_9938_), .B(_9939_), .Y(_9940_) );
	NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_9940_), .Y(_9941_) );
	OAI21X1 OAI21X1_4155 ( .gnd(gnd), .vdd(vdd), .A(_9941_), .B(_9700_), .C(csr_gpr_iu_csr_mtvec_24_), .Y(_9942_) );
	NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_9941_), .B(_9700_), .Y(_9943_) );
	NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9943_), .Y(_9944_) );
	AOI21X1 AOI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_9944_), .B(_9942_), .C(_9275_), .Y(_9945_) );
	OAI22X1 OAI22X1_769 ( .gnd(gnd), .vdd(vdd), .A(_9073_), .B(_9280_), .C(_9925_), .D(_9274_), .Y(_9946_) );
	OAI21X1 OAI21X1_4156 ( .gnd(gnd), .vdd(vdd), .A(_9946_), .B(_9945_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf1), .Y(_9947_) );
	NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_9917_), .B(_9913_), .Y(_9948_) );
	OAI21X1 OAI21X1_4157 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_24_), .B(_9914_), .C(_9322__bF_buf3), .Y(_9949_) );
	OAI21X1 OAI21X1_4158 ( .gnd(gnd), .vdd(vdd), .A(_9917_), .B(_9285__bF_buf3), .C(_9149__bF_buf4), .Y(_9950_) );
	AOI21X1 AOI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_25_), .B(_9326_), .C(_9950_), .Y(_9951_) );
	OAI21X1 OAI21X1_4159 ( .gnd(gnd), .vdd(vdd), .A(_9948_), .B(_9949_), .C(_9951_), .Y(_9952_) );
	OAI21X1 OAI21X1_4160 ( .gnd(gnd), .vdd(vdd), .A(_7424__bF_buf2), .B(_8615_), .C(_9952_), .Y(_9953_) );
	OAI21X1 OAI21X1_4161 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .B(_9149__bF_buf3), .C(_9251__bF_buf4), .Y(_9954_) );
	AOI21X1 AOI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_9953_), .B(_9947_), .C(_9954_), .Y(_9955_) );
	OAI21X1 OAI21X1_4162 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9251__bF_buf3), .C(_9095__bF_buf1), .Y(_9956_) );
	NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .B(_9097_), .Y(_9957_) );
	OAI21X1 OAI21X1_4163 ( .gnd(gnd), .vdd(vdd), .A(_8977_), .B(_9105__bF_buf3), .C(_9957_), .Y(_9958_) );
	AOI21X1 AOI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_24_), .B(_9098__bF_buf3), .C(_9958_), .Y(_9959_) );
	AOI21X1 AOI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_9959_), .B(_9094__bF_buf1), .C(_7303__bF_buf12_bF_buf3), .Y(_9960_) );
	OAI21X1 OAI21X1_4164 ( .gnd(gnd), .vdd(vdd), .A(_9956_), .B(_9955_), .C(_9960_), .Y(_9961_) );
	AOI21X1 AOI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_9937_), .B(_9961_), .C(rst_bF_buf23), .Y(_6725__24_) );
	INVX1 INVX1_1667 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_25_), .Y(_9962_) );
	AOI21X1 AOI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf5), .B(_9962_), .C(_7304__bF_buf10_bF_buf3), .Y(_9963_) );
	OAI21X1 OAI21X1_4165 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .B(_9268__bF_buf4), .C(_9963_), .Y(_9964_) );
	OAI21X1 OAI21X1_4166 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_31_), .B(csr_gpr_iu_csr_mtvec_26_), .C(_9274_), .Y(_9965_) );
	INVX1 INVX1_1668 ( .gnd(gnd), .vdd(vdd), .A(_9965_), .Y(_9966_) );
	AOI21X1 AOI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_9501_), .B(_9502_), .C(_9698_), .Y(_9967_) );
	NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_9697_), .B(_9695_), .Y(_9968_) );
	INVX1 INVX1_1669 ( .gnd(gnd), .vdd(vdd), .A(_9968_), .Y(_9969_) );
	INVX1 INVX1_1670 ( .gnd(gnd), .vdd(vdd), .A(_9941_), .Y(_9970_) );
	OAI21X1 OAI21X1_4167 ( .gnd(gnd), .vdd(vdd), .A(_9967_), .B(_9969_), .C(_9970_), .Y(_9971_) );
	OAI21X1 OAI21X1_4168 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9971_), .C(csr_gpr_iu_csr_mtvec_25_), .Y(_9972_) );
	NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_24_), .B(_9073_), .C(_9943_), .Y(_9973_) );
	NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_31_), .B(_9972_), .C(_9973_), .Y(_9974_) );
	AOI22X1 AOI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_25_), .B(_9273__bF_buf0), .C(_9966_), .D(_9974_), .Y(_9975_) );
	NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_25_), .B(_9948_), .Y(_9976_) );
	NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_9917_), .B(_8095_), .Y(_9977_) );
	INVX1 INVX1_1671 ( .gnd(gnd), .vdd(vdd), .A(_9977_), .Y(_9978_) );
	OAI21X1 OAI21X1_4169 ( .gnd(gnd), .vdd(vdd), .A(_9978_), .B(_9913_), .C(_9322__bF_buf2), .Y(_9979_) );
	OAI21X1 OAI21X1_4170 ( .gnd(gnd), .vdd(vdd), .A(_8095_), .B(_9285__bF_buf2), .C(_9149__bF_buf2), .Y(_9980_) );
	AOI21X1 AOI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_26_), .B(_9326_), .C(_9980_), .Y(_9981_) );
	OAI21X1 OAI21X1_4171 ( .gnd(gnd), .vdd(vdd), .A(_9979_), .B(_9976_), .C(_9981_), .Y(_9982_) );
	OAI21X1 OAI21X1_4172 ( .gnd(gnd), .vdd(vdd), .A(_7424__bF_buf1), .B(_8615_), .C(_9982_), .Y(_9983_) );
	OAI21X1 OAI21X1_4173 ( .gnd(gnd), .vdd(vdd), .A(_8613_), .B(_9975_), .C(_9983_), .Y(_9984_) );
	AOI21X1 AOI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_7875_), .C(_9292_), .Y(_9985_) );
	OAI21X1 OAI21X1_4174 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .B(_9251__bF_buf2), .C(_9095__bF_buf0), .Y(_9986_) );
	AOI21X1 AOI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_9984_), .B(_9985_), .C(_9986_), .Y(_9987_) );
	NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf3), .B(_9103_), .Y(_9988_) );
	AOI22X1 AOI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .B(_9097_), .C(csr_gpr_iu_csr_mepc_25_), .D(_9104_), .Y(_9989_) );
	OAI21X1 OAI21X1_4175 ( .gnd(gnd), .vdd(vdd), .A(_7872_), .B(_9988_), .C(_9989_), .Y(_9990_) );
	OAI21X1 OAI21X1_4176 ( .gnd(gnd), .vdd(vdd), .A(_9990_), .B(_9095__bF_buf4), .C(_7304__bF_buf9_bF_buf3), .Y(_9991_) );
	OAI21X1 OAI21X1_4177 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .B(_9987_), .C(_9964_), .Y(_9992_) );
	AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_9992_), .B(_6879__bF_buf13), .Y(_6725__25_) );
	INVX1 INVX1_1672 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_26_), .Y(_9993_) );
	AOI21X1 AOI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf3), .B(_9993_), .C(_7304__bF_buf8_bF_buf3), .Y(_9994_) );
	OAI21X1 OAI21X1_4178 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(_9268__bF_buf2), .C(_9994_), .Y(_9995_) );
	AOI21X1 AOI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_9914_), .B(_9977_), .C(csr_gpr_iu_csr_stvec_26_), .Y(_9996_) );
	NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_26_), .B(_9977_), .Y(_9997_) );
	OAI21X1 OAI21X1_4179 ( .gnd(gnd), .vdd(vdd), .A(_9997_), .B(_9913_), .C(_9322__bF_buf1), .Y(_9998_) );
	INVX1 INVX1_1673 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_26_), .Y(_9999_) );
	OAI21X1 OAI21X1_4180 ( .gnd(gnd), .vdd(vdd), .A(_9999_), .B(_9285__bF_buf1), .C(_9149__bF_buf1), .Y(_10000_) );
	AOI21X1 AOI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_27_), .B(_9326_), .C(_10000_), .Y(_10001_) );
	OAI21X1 OAI21X1_4181 ( .gnd(gnd), .vdd(vdd), .A(_9998_), .B(_9996_), .C(_10001_), .Y(_10002_) );
	OAI21X1 OAI21X1_4182 ( .gnd(gnd), .vdd(vdd), .A(_8613_), .B(_9291_), .C(_10002_), .Y(_10003_) );
	NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9073_), .Y(_10004_) );
	AOI21X1 AOI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_10004_), .C(csr_gpr_iu_csr_mtvec_26_), .Y(_10005_) );
	NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_26_), .B(_10004_), .C(_9943_), .Y(_10006_) );
	NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_9276__bF_buf1), .B(_10006_), .Y(_10007_) );
	NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_10005_), .B(_10007_), .Y(_10008_) );
	NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_26_), .B(_9273__bF_buf3), .Y(_10009_) );
	OAI21X1 OAI21X1_4183 ( .gnd(gnd), .vdd(vdd), .A(_9077_), .B(_9280_), .C(_10009_), .Y(_10010_) );
	OAI21X1 OAI21X1_4184 ( .gnd(gnd), .vdd(vdd), .A(_10010_), .B(_10008_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf0), .Y(_10011_) );
	OAI21X1 OAI21X1_4185 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(_9149__bF_buf0), .C(_9251__bF_buf1), .Y(_10012_) );
	AOI21X1 AOI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_10011_), .B(_10003_), .C(_10012_), .Y(_10013_) );
	OAI21X1 OAI21X1_4186 ( .gnd(gnd), .vdd(vdd), .A(_9993_), .B(_9251__bF_buf0), .C(_9095__bF_buf3), .Y(_10014_) );
	NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_26_), .B(_9098__bF_buf2), .Y(_10015_) );
	OAI21X1 OAI21X1_4187 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(biu_mmu_msu_0_bF_buf2), .C(_10015_), .Y(_10016_) );
	AOI21X1 AOI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_26_), .B(_9104_), .C(_10016_), .Y(_10017_) );
	AOI21X1 AOI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf0), .B(_10017_), .C(_7303__bF_buf11_bF_buf3), .Y(_10018_) );
	OAI21X1 OAI21X1_4188 ( .gnd(gnd), .vdd(vdd), .A(_10014_), .B(_10013_), .C(_10018_), .Y(_10019_) );
	AOI21X1 AOI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_10019_), .B(_9995_), .C(rst_bF_buf22), .Y(_6725__26_) );
	INVX1 INVX1_1674 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_27_), .Y(_10020_) );
	AOI21X1 AOI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf1), .B(_10020_), .C(_7304__bF_buf7_bF_buf3), .Y(_10021_) );
	OAI21X1 OAI21X1_4189 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .B(_9268__bF_buf0), .C(_10021_), .Y(_10022_) );
	OAI21X1 OAI21X1_4190 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_9285__bF_buf0), .C(_9149__bF_buf4), .Y(_10023_) );
	NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_9997_), .B(_9913_), .Y(_10024_) );
	NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_26_), .B(csr_gpr_iu_csr_stvec_27_), .Y(_10025_) );
	NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_10025_), .B(_9978_), .Y(_10026_) );
	NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_9912_), .B(_10026_), .C(_9759_), .Y(_10027_) );
	OAI21X1 OAI21X1_4191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_27_), .B(_10024_), .C(_10027_), .Y(_10028_) );
	OAI21X1 OAI21X1_4192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf2), .B(csr_gpr_iu_csr_stvec_28_), .C(_9285__bF_buf4), .Y(_10029_) );
	AOI21X1 AOI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_10028_), .B(csr_gpr_iu_csr_scause_31_bF_buf1), .C(_10029_), .Y(_10030_) );
	OAI21X1 OAI21X1_4193 ( .gnd(gnd), .vdd(vdd), .A(_10023_), .B(_10030_), .C(_8861__bF_buf1), .Y(_10031_) );
	INVX1 INVX1_1675 ( .gnd(gnd), .vdd(vdd), .A(_10004_), .Y(_10032_) );
	NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_26_), .B(csr_gpr_iu_csr_mtvec_27_), .Y(_10033_) );
	NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_10033_), .B(_10032_), .Y(_10034_) );
	INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(_10034_), .Y(_10035_) );
	OAI21X1 OAI21X1_4194 ( .gnd(gnd), .vdd(vdd), .A(_10035_), .B(_9971_), .C(_9276__bF_buf0), .Y(_10036_) );
	AOI21X1 AOI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_10006_), .B(_9077_), .C(_10036_), .Y(_10037_) );
	INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_28_), .Y(_10038_) );
	OAI22X1 OAI22X1_770 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9280_), .C(_9077_), .D(_9274_), .Y(_10039_) );
	OAI21X1 OAI21X1_4195 ( .gnd(gnd), .vdd(vdd), .A(_10039_), .B(_10037_), .C(csr_gpr_iu_csr_priv_d_1_bF_buf3), .Y(_10040_) );
	OAI21X1 OAI21X1_4196 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .B(_9149__bF_buf3), .C(_9251__bF_buf6), .Y(_10041_) );
	AOI21X1 AOI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_10031_), .B(_10040_), .C(_10041_), .Y(_10042_) );
	OAI21X1 OAI21X1_4197 ( .gnd(gnd), .vdd(vdd), .A(_10020_), .B(_9251__bF_buf5), .C(_9095__bF_buf2), .Y(_10043_) );
	NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .B(_9097_), .Y(_10044_) );
	OAI21X1 OAI21X1_4198 ( .gnd(gnd), .vdd(vdd), .A(_7895_), .B(_9988_), .C(_10044_), .Y(_10045_) );
	AOI21X1 AOI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_27_), .B(_9104_), .C(_10045_), .Y(_10046_) );
	AOI21X1 AOI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf5), .B(_10046_), .C(_7303__bF_buf10_bF_buf3), .Y(_10047_) );
	OAI21X1 OAI21X1_4199 ( .gnd(gnd), .vdd(vdd), .A(_10043_), .B(_10042_), .C(_10047_), .Y(_10048_) );
	AOI21X1 AOI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_10048_), .B(_10022_), .C(rst_bF_buf21), .Y(_6725__27_) );
	INVX1 INVX1_1676 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .Y(_10049_) );
	OAI21X1 OAI21X1_4200 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9246_), .C(csr_gpr_iu_csr_pc_next_28_), .Y(_10050_) );
	OAI21X1 OAI21X1_4201 ( .gnd(gnd), .vdd(vdd), .A(_10049_), .B(_9268__bF_buf6), .C(_10050_), .Y(_10051_) );
	NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf9_bF_buf3), .B(_10051_), .Y(_10052_) );
	INVX1 INVX1_1677 ( .gnd(gnd), .vdd(vdd), .A(_10026_), .Y(_10053_) );
	NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_9911_), .B(_10053_), .C(_9713_), .Y(_10054_) );
	NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_28_), .B(_10054_), .Y(_10055_) );
	INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_28_), .Y(_10056_) );
	NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_27_), .B(_10024_), .Y(_10057_) );
	OAI21X1 OAI21X1_4202 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_10057_), .C(_9322__bF_buf0), .Y(_10058_) );
	OAI21X1 OAI21X1_4203 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_9285__bF_buf3), .C(_9149__bF_buf2), .Y(_10059_) );
	AOI21X1 AOI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_29_), .B(_9326_), .C(_10059_), .Y(_10060_) );
	OAI21X1 OAI21X1_4204 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .B(_10058_), .C(_10060_), .Y(_10061_) );
	OAI21X1 OAI21X1_4205 ( .gnd(gnd), .vdd(vdd), .A(_10035_), .B(_9971_), .C(_10038_), .Y(_10062_) );
	NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_10035_), .B(_9971_), .Y(_10063_) );
	NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_28_), .B(_10063_), .Y(_10064_) );
	NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_10062_), .B(_10064_), .Y(_10065_) );
	AOI22X1 AOI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_28_), .B(_9273__bF_buf2), .C(csr_gpr_iu_csr_mtvec_29_), .D(_9281__bF_buf1), .Y(_10066_) );
	OAI21X1 OAI21X1_4206 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_10065_), .C(_10066_), .Y(_10067_) );
	AOI22X1 AOI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(_10061_), .B(_8861__bF_buf0), .C(csr_gpr_iu_csr_priv_d_1_bF_buf2), .D(_10067_), .Y(_10068_) );
	OAI21X1 OAI21X1_4207 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .B(_9149__bF_buf1), .C(_9251__bF_buf4), .Y(_10069_) );
	AOI21X1 AOI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(csr_gpr_iu_csr_pc_next_28_), .C(_9094__bF_buf4), .Y(_10070_) );
	OAI21X1 OAI21X1_4208 ( .gnd(gnd), .vdd(vdd), .A(_10069_), .B(_10068_), .C(_10070_), .Y(_10071_) );
	OAI22X1 OAI22X1_771 ( .gnd(gnd), .vdd(vdd), .A(_10049_), .B(biu_mmu_msu_0_bF_buf1), .C(_7904_), .D(_9988_), .Y(_10072_) );
	AOI21X1 AOI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_28_), .B(_9104_), .C(_10072_), .Y(_10073_) );
	AOI21X1 AOI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf3), .B(_10073_), .C(_7303__bF_buf8_bF_buf3), .Y(_10074_) );
	NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_10074_), .B(_10071_), .Y(_10075_) );
	AOI21X1 AOI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_10075_), .B(_10052_), .C(rst_bF_buf20), .Y(_6725__28_) );
	INVX1 INVX1_1678 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_29_), .Y(_10076_) );
	AOI21X1 AOI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_9268__bF_buf5), .B(_10076_), .C(_7304__bF_buf6_bF_buf3), .Y(_10077_) );
	OAI21X1 OAI21X1_4209 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(_9268__bF_buf4), .C(_10077_), .Y(_10078_) );
	AOI21X1 AOI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_10063_), .B(csr_gpr_iu_csr_mtvec_28_), .C(csr_gpr_iu_csr_mtvec_29_), .Y(_10079_) );
	OAI21X1 OAI21X1_4210 ( .gnd(gnd), .vdd(vdd), .A(_9081_), .B(_10064_), .C(_9276__bF_buf3), .Y(_10080_) );
	AOI22X1 AOI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_29_), .B(_9273__bF_buf1), .C(csr_gpr_iu_csr_mtvec_30_), .D(_9281__bF_buf0), .Y(_10081_) );
	OAI21X1 OAI21X1_4211 ( .gnd(gnd), .vdd(vdd), .A(_10079_), .B(_10080_), .C(_10081_), .Y(_10082_) );
	NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_10082_), .Y(_10083_) );
	OAI21X1 OAI21X1_4212 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_priv_d_0_), .B(_7936_), .C(_7427_), .Y(_10084_) );
	AOI21X1 AOI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_29_), .B(_9284_), .C(_7427_), .Y(_10085_) );
	OAI21X1 OAI21X1_4213 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_10027_), .C(_8101_), .Y(_10086_) );
	NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_28_), .B(csr_gpr_iu_csr_stvec_29_), .C(_10054_), .Y(_10087_) );
	AOI21X1 AOI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_10087_), .B(_10086_), .C(_7571_), .Y(_10088_) );
	OAI21X1 OAI21X1_4214 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf0), .B(csr_gpr_iu_csr_stvec_30_), .C(_9285__bF_buf2), .Y(_10089_) );
	OAI21X1 OAI21X1_4215 ( .gnd(gnd), .vdd(vdd), .A(_10089_), .B(_10088_), .C(_10085_), .Y(_10090_) );
	AOI21X1 AOI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_10090_), .B(_10084_), .C(_7424__bF_buf0), .Y(_10091_) );
	OAI21X1 OAI21X1_4216 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(_7423_), .C(_9251__bF_buf3), .Y(_10092_) );
	AOI21X1 AOI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_10091_), .B(_10083_), .C(_10092_), .Y(_10093_) );
	OAI21X1 OAI21X1_4217 ( .gnd(gnd), .vdd(vdd), .A(_10076_), .B(_9251__bF_buf2), .C(_9095__bF_buf1), .Y(_10094_) );
	OAI22X1 OAI22X1_772 ( .gnd(gnd), .vdd(vdd), .A(_7936_), .B(biu_mmu_msu_0_bF_buf0), .C(_7913_), .D(_9988_), .Y(_10095_) );
	AOI21X1 AOI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_29_), .B(_9104_), .C(_10095_), .Y(_10096_) );
	AOI21X1 AOI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf2), .B(_10096_), .C(_7303__bF_buf7_bF_buf3), .Y(_10097_) );
	OAI21X1 OAI21X1_4218 ( .gnd(gnd), .vdd(vdd), .A(_10094_), .B(_10093_), .C(_10097_), .Y(_10098_) );
	AOI21X1 AOI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_10098_), .B(_10078_), .C(rst_bF_buf19), .Y(_6725__29_) );
	OAI21X1 OAI21X1_4219 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9246_), .C(csr_gpr_iu_csr_pc_next_30_), .Y(_10099_) );
	OAI21X1 OAI21X1_4220 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(_9268__bF_buf3), .C(_10099_), .Y(_10100_) );
	NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_7303__bF_buf6_bF_buf3), .B(_10100_), .Y(_10101_) );
	INVX1 INVX1_1679 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_30_), .Y(_10102_) );
	NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9081_), .Y(_10103_) );
	AOI21X1 AOI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_10063_), .B(_10103_), .C(_10102_), .Y(_10104_) );
	NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_10034_), .B(_10103_), .C(_9943_), .Y(_10105_) );
	NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_30_), .B(_10105_), .Y(_10106_) );
	OAI21X1 OAI21X1_4221 ( .gnd(gnd), .vdd(vdd), .A(_10106_), .B(_10104_), .C(_9276__bF_buf2), .Y(_10107_) );
	AOI22X1 AOI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_30_), .B(_9273__bF_buf0), .C(csr_gpr_iu_csr_mtvec_31_), .D(_9281__bF_buf3), .Y(_10108_) );
	AOI21X1 AOI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_10107_), .B(_10108_), .C(_8615_), .Y(_10109_) );
	OAI21X1 OAI21X1_4222 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(_7426_), .C(_8615_), .Y(_10110_) );
	INVX1 INVX1_1680 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_30_), .Y(_10111_) );
	OAI21X1 OAI21X1_4223 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_9285__bF_buf1), .C(_7426_), .Y(_10112_) );
	NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_8101_), .Y(_10113_) );
	INVX1 INVX1_1681 ( .gnd(gnd), .vdd(vdd), .A(_10113_), .Y(_10114_) );
	OAI21X1 OAI21X1_4224 ( .gnd(gnd), .vdd(vdd), .A(_10114_), .B(_10027_), .C(csr_gpr_iu_csr_stvec_30_), .Y(_10115_) );
	NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10113_), .C(_10054_), .Y(_10116_) );
	NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf3), .B(_10115_), .C(_10116_), .Y(_10117_) );
	OAI21X1 OAI21X1_4225 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_31_bF_buf2), .B(csr_gpr_iu_csr_stvec_31_), .C(_9285__bF_buf0), .Y(_10118_) );
	INVX1 INVX1_1682 ( .gnd(gnd), .vdd(vdd), .A(_10118_), .Y(_10119_) );
	AOI21X1 AOI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_10117_), .B(_10119_), .C(_10112_), .Y(_10120_) );
	OAI21X1 OAI21X1_4226 ( .gnd(gnd), .vdd(vdd), .A(_10110_), .B(_10120_), .C(_7423_), .Y(_10121_) );
	AOI21X1 AOI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(_7424__bF_buf3), .C(_9292_), .Y(_10122_) );
	OAI21X1 OAI21X1_4227 ( .gnd(gnd), .vdd(vdd), .A(_10109_), .B(_10121_), .C(_10122_), .Y(_10123_) );
	AOI21X1 AOI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(csr_gpr_iu_csr_pc_next_30_), .C(_9094__bF_buf1), .Y(_10124_) );
	NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_10123_), .Y(_10125_) );
	OAI22X1 OAI22X1_773 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(biu_mmu_msu_0_bF_buf4), .C(_7935_), .D(_9988_), .Y(_10126_) );
	AOI21X1 AOI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_30_), .B(_9104_), .C(_10126_), .Y(_10127_) );
	AOI21X1 AOI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf0), .B(_10127_), .C(_7303__bF_buf5_bF_buf3), .Y(_10128_) );
	NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_10128_), .B(_10125_), .Y(_10129_) );
	AOI21X1 AOI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_10129_), .B(_10101_), .C(rst_bF_buf18), .Y(_6725__30_) );
	INVX1 INVX1_1683 ( .gnd(gnd), .vdd(vdd), .A(_10103_), .Y(_10130_) );
	NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_10035_), .B(_10130_), .C(_9971_), .Y(_10131_) );
	AOI21X1 AOI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_10131_), .B(csr_gpr_iu_csr_mtvec_30_), .C(_9085_), .Y(_10132_) );
	NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_10102_), .B(csr_gpr_iu_csr_mtvec_31_), .C(_10105_), .Y(_10133_) );
	OAI21X1 OAI21X1_4228 ( .gnd(gnd), .vdd(vdd), .A(_10133_), .B(_10132_), .C(_9276__bF_buf1), .Y(_10134_) );
	NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_31_), .B(_9273__bF_buf3), .Y(_10135_) );
	NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_10135_), .C(_10134_), .Y(_10136_) );
	NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_10114_), .B(_10027_), .Y(_10137_) );
	AOI21X1 AOI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_10137_), .B(csr_gpr_iu_csr_stvec_30_), .C(_8104_), .Y(_10138_) );
	NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_10113_), .B(_10054_), .Y(_10139_) );
	NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(csr_gpr_iu_csr_stvec_31_), .C(_10139_), .Y(_10140_) );
	OAI21X1 OAI21X1_4229 ( .gnd(gnd), .vdd(vdd), .A(_10138_), .B(_10140_), .C(_9322__bF_buf3), .Y(_10141_) );
	NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_31_), .B(_9284_), .Y(_10142_) );
	NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_7426_), .B(_10142_), .C(_10141_), .Y(_10143_) );
	INVX1 INVX1_1684 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .Y(_10144_) );
	AOI21X1 AOI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_10144_), .C(_7424__bF_buf2), .Y(_10145_) );
	NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_10145_), .B(_10136_), .C(_10143_), .Y(_10146_) );
	AOI21X1 AOI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .B(_7424__bF_buf1), .C(_9292_), .Y(_10147_) );
	NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_10147_), .B(_10146_), .Y(_10148_) );
	INVX1 INVX1_1685 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_31_), .Y(_10149_) );
	AOI21X1 AOI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_10149_), .C(_9094__bF_buf5), .Y(_10150_) );
	NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_10150_), .B(_10148_), .Y(_10151_) );
	OAI22X1 OAI22X1_774 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .B(biu_mmu_msu_0_bF_buf3), .C(csr_gpr_iu_csr_sepc_31_), .D(_9988_), .Y(_10152_) );
	AOI21X1 AOI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_9014_), .B(_9104_), .C(_10152_), .Y(_10153_) );
	AOI21X1 AOI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_9094__bF_buf4), .B(_10153_), .C(_7303__bF_buf4_bF_buf3), .Y(_10154_) );
	NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9247_), .Y(_10155_) );
	OAI21X1 OAI21X1_4230 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9268__bF_buf2), .C(_7303__bF_buf3_bF_buf3), .Y(_10156_) );
	OAI21X1 OAI21X1_4231 ( .gnd(gnd), .vdd(vdd), .A(_10155_), .B(_10156_), .C(_6879__bF_buf12), .Y(_10157_) );
	AOI21X1 AOI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_10151_), .B(_10154_), .C(_10157_), .Y(_6725__31_) );
	NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(_6813_), .Y(_10158_) );
	NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_10158_), .B(_8109_), .Y(_10159_) );
	INVX1 INVX1_1686 ( .gnd(gnd), .vdd(vdd), .A(_10159_), .Y(_10160_) );
	NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_8057_), .B(_10160_), .Y(_10161_) );
	NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_10161_), .Y(_10162_) );
	INVX8 INVX8_88 ( .gnd(gnd), .vdd(vdd), .A(_9019__bF_buf0), .Y(_10163_) );
	NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_7313_), .B(_10161_), .Y(_10164_) );
	INVX4 INVX4_26 ( .gnd(gnd), .vdd(vdd), .A(_10164_), .Y(_10165_) );
	AOI22X1 AOI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_0_), .B(_10163_), .C(csr_gpr_iu_csr_mcycle_0_), .D(_10165_), .Y(_10166_) );
	OAI21X1 OAI21X1_4232 ( .gnd(gnd), .vdd(vdd), .A(_6822_), .B(_10162_), .C(_10166_), .Y(_10167_) );
	AOI22X1 AOI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf2), .B(biu_mmu_ag0_12_), .C(csr_gpr_iu_csr_stvec_0_), .D(_8062__bF_buf5), .Y(_10168_) );
	OAI21X1 OAI21X1_4233 ( .gnd(gnd), .vdd(vdd), .A(_8685_), .B(_8684__bF_buf3), .C(_10168_), .Y(_10169_) );
	INVX4 INVX4_27 ( .gnd(gnd), .vdd(vdd), .A(_8486__bF_buf0), .Y(_10170_) );
	OAI21X1 OAI21X1_4234 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_0_), .B(csr_gpr_iu_csr_mideleg_0_), .C(_10170_), .Y(_10171_) );
	OAI21X1 OAI21X1_4235 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_7959_), .C(_10171_), .Y(_10172_) );
	OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_10172_), .B(_10169_), .Y(_10173_) );
	NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_10167_), .B(_10173_), .Y(_10174_) );
	AOI22X1 AOI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf3), .B(csr_gpr_iu_csr_sscratch_0_), .C(csr_gpr_iu_csr_sepc_0_), .D(_7584__bF_buf0), .Y(_10175_) );
	AOI22X1 AOI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_0_), .B(_8417__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr0_0_), .D(_8280__bF_buf0), .Y(_10176_) );
	AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_10175_), .Y(_10177_) );
	AOI22X1 AOI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_0_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_mtval_0_), .D(_8618__bF_buf2), .Y(_10178_) );
	AOI22X1 AOI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_0_), .B(_8846__bF_buf0), .C(csr_gpr_iu_csr_pmp0cfg_0_), .D(_8372__bF_buf4), .Y(_10179_) );
	NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_10179_), .B(_10178_), .Y(_10180_) );
	AOI22X1 AOI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_0_), .B(_7435__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_0_), .D(_8117__bF_buf4), .Y(_10181_) );
	INVX8 INVX8_89 ( .gnd(gnd), .vdd(vdd), .A(_8162__bF_buf2), .Y(_10182_) );
	AOI22X1 AOI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp4cfg_0_), .B(_8327__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr2_0_), .D(_10182__bF_buf3), .Y(_10183_) );
	NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_10181_), .B(_10183_), .Y(_10184_) );
	NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_10180_), .B(_10184_), .Y(_10185_) );
	NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_10177_), .B(_10185_), .C(_10174_), .Y(csr_0_) );
	NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_10160_), .Y(_10186_) );
	AOI22X1 AOI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf3), .B(csr_gpr_iu_csr_sie), .C(csr_gpr_iu_csr_mcycle_1_), .D(_10186_), .Y(_10187_) );
	NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_1_), .B(_10163_), .Y(_10188_) );
	NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_1_), .B(_8417__bF_buf4), .Y(_10189_) );
	AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10188_), .Y(_10190_) );
	AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_10190_), .B(_10187_), .Y(_10191_) );
	NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_1_), .B(_8117__bF_buf3), .Y(_10192_) );
	AOI22X1 AOI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_ssie), .B(_8469_), .C(csr_gpr_iu_csr_sie), .D(_9144_), .Y(_10193_) );
	NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_10193_), .B(_10192_), .Y(_10194_) );
	NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_8466_), .B(_8845_), .Y(_10195_) );
	NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .B(_10195_), .Y(_10196_) );
	NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_8106_), .Y(_10197_) );
	NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .B(_10197_), .Y(_10198_) );
	INVX4 INVX4_28 ( .gnd(gnd), .vdd(vdd), .A(_10198_), .Y(_10199_) );
	AOI22X1 AOI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_13_), .B(_9234__bF_buf1), .C(csr_gpr_iu_csr_stval_1_), .D(_10199_), .Y(_10200_) );
	OAI21X1 OAI21X1_4236 ( .gnd(gnd), .vdd(vdd), .A(_7284_), .B(_10196_), .C(_10200_), .Y(_10201_) );
	OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_10194_), .B(_10201_), .Y(_10202_) );
	NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_1_), .B(_8062__bF_buf4), .Y(_10203_) );
	AOI22X1 AOI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_1_), .B(_8165__bF_buf1), .C(csr_gpr_iu_csr_scause_1_), .D(_7435__bF_buf0), .Y(_10204_) );
	AOI22X1 AOI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf2), .B(csr_gpr_iu_csr_sscratch_1_), .C(csr_gpr_iu_csr_sepc_1_), .D(_7584__bF_buf5), .Y(_10205_) );
	NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_10203_), .B(_10204_), .C(_10205_), .Y(_10206_) );
	NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_10206_), .B(_10202_), .Y(_10207_) );
	NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_10160_), .B(_8488_), .Y(_10208_) );
	INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(_10208_), .Y(_10209_) );
	AOI22X1 AOI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp0cfg_1_), .B(_8372__bF_buf3), .C(csr_gpr_iu_csr_pmp4cfg_1_), .D(_8327__bF_buf3), .Y(_10210_) );
	OAI21X1 OAI21X1_4237 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_1_), .B(csr_gpr_iu_csr_mideleg_1_), .C(_8489__bF_buf0), .Y(_10211_) );
	AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_10210_), .B(_10211_), .Y(_10212_) );
	OAI21X1 OAI21X1_4238 ( .gnd(gnd), .vdd(vdd), .A(_6881_), .B(_10209_), .C(_10212_), .Y(_10213_) );
	NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf2), .B(_7434__bF_buf1), .Y(_10214_) );
	INVX4 INVX4_29 ( .gnd(gnd), .vdd(vdd), .A(_10214_), .Y(_10215_) );
	OAI22X1 OAI22X1_775 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .B(_8847__bF_buf7), .C(_8690_), .D(_10215_), .Y(_10216_) );
	AOI21X1 AOI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_1_), .B(_8233__bF_buf0), .C(_10216_), .Y(_10217_) );
	NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .B(_10195_), .Y(_10218_) );
	OAI22X1 OAI22X1_776 ( .gnd(gnd), .vdd(vdd), .A(_7284_), .B(_10218_), .C(_8622_), .D(_8617_), .Y(_10219_) );
	AOI21X1 AOI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_1_), .B(_8280__bF_buf5), .C(_10219_), .Y(_10220_) );
	NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_10220_), .B(_10217_), .Y(_10221_) );
	NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .B(_10213_), .Y(_10222_) );
	NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_10191_), .B(_10207_), .C(_10222_), .Y(csr_1_) );
	INVX1 INVX1_1687 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_14_), .Y(_10223_) );
	AOI22X1 AOI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_2_), .B(_8062__bF_buf3), .C(csr_gpr_iu_csr_mcycle_2_), .D(_10165_), .Y(_10224_) );
	OAI21X1 OAI21X1_4239 ( .gnd(gnd), .vdd(vdd), .A(_10223_), .B(_9161__bF_buf4), .C(_10224_), .Y(_10225_) );
	OAI21X1 OAI21X1_4240 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_2_), .B(csr_gpr_iu_csr_mideleg_2_), .C(_10170_), .Y(_10226_) );
	INVX4 INVX4_30 ( .gnd(gnd), .vdd(vdd), .A(_10162_), .Y(_10227_) );
	AOI22X1 AOI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_2_), .B(_10163_), .C(csr_gpr_iu_csr_minstret_2_), .D(_10227_), .Y(_10228_) );
	AOI22X1 AOI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr2_2_), .C(csr_gpr_iu_csr_mtval_2_), .D(_8618__bF_buf1), .Y(_10229_) );
	NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_10226_), .B(_10229_), .C(_10228_), .Y(_10230_) );
	NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_10225_), .B(_10230_), .Y(_10231_) );
	AOI22X1 AOI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_2_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_stval_2_), .D(_7960__bF_buf3), .Y(_10232_) );
	AOI22X1 AOI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp4cfg_2_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmp0cfg_2_), .D(_8372__bF_buf2), .Y(_10233_) );
	AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_10232_), .B(_10233_), .Y(_10234_) );
	INVX4 INVX4_31 ( .gnd(gnd), .vdd(vdd), .A(_8684__bF_buf2), .Y(_10235_) );
	AOI22X1 AOI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf4), .B(csr_gpr_iu_csr_sepc_2_), .C(csr_gpr_iu_csr_mcause_2_), .D(_10235_), .Y(_10236_) );
	AOI22X1 AOI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf6), .B(csr_gpr_iu_csr_scause_2_), .C(csr_gpr_iu_csr_pmpaddr1_2_), .D(_8233__bF_buf5), .Y(_10237_) );
	NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_10237_), .B(_10236_), .Y(_10238_) );
	AOI22X1 AOI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_2_), .B(_8846__bF_buf3), .C(csr_gpr_iu_csr_mscratch_2_), .D(_8417__bF_buf3), .Y(_10239_) );
	AOI22X1 AOI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_2_), .B(_7323__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr0_2_), .D(_8280__bF_buf4), .Y(_10240_) );
	NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_10239_), .B(_10240_), .Y(_10241_) );
	NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_10238_), .B(_10241_), .Y(_10242_) );
	NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_10234_), .B(_10242_), .C(_10231_), .Y(csr_2_) );
	INVX1 INVX1_1688 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp4cfg_3_), .Y(_10243_) );
	NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_8111__bF_buf1), .B(_8468_), .Y(_10244_) );
	AOI22X1 AOI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_msie), .B(_10244_), .C(csr_gpr_iu_csr_mscratch_3_), .D(_8417__bF_buf2), .Y(_10245_) );
	OAI21X1 OAI21X1_4241 ( .gnd(gnd), .vdd(vdd), .A(_9028_), .B(_9019__bF_buf5), .C(_10245_), .Y(_10246_) );
	NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_3_), .B(_10208_), .Y(_10247_) );
	OAI21X1 OAI21X1_4242 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_3_), .B(csr_gpr_iu_csr_mideleg_3_), .C(_8489__bF_buf5), .Y(_10248_) );
	AOI22X1 AOI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf2), .B(csr_gpr_iu_csr_mie), .C(csr_gpr_iu_csr_mcycle_3_), .D(_10186_), .Y(_10249_) );
	NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(_10247_), .C(_10248_), .Y(_10250_) );
	NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_10250_), .B(_10246_), .Y(_10251_) );
	OAI21X1 OAI21X1_4243 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .B(_8326_), .C(_10251_), .Y(_10252_) );
	AOI22X1 AOI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_15_), .B(_9234__bF_buf0), .C(csr_gpr_iu_csr_stval_3_), .D(_10199_), .Y(_10253_) );
	AOI22X1 AOI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf3), .B(csr_gpr_iu_csr_sepc_3_), .C(csr_gpr_iu_csr_scause_3_), .D(_7435__bF_buf5), .Y(_10254_) );
	NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_10254_), .B(_10253_), .Y(_10255_) );
	AOI22X1 AOI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_3_), .B(_7319__bF_buf1), .C(csr_gpr_iu_csr_stvec_3_), .D(_8062__bF_buf2), .Y(_10256_) );
	AOI22X1 AOI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(_8117__bF_buf1), .B(csr_gpr_iu_csr_pmpaddr3_3_), .C(csr_gpr_iu_csr_pmpaddr2_3_), .D(_10182__bF_buf1), .Y(_10257_) );
	NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_10256_), .B(_10257_), .Y(_10258_) );
	NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_10258_), .Y(_10259_) );
	AOI22X1 AOI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_3_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr0_3_), .D(_8280__bF_buf3), .Y(_10260_) );
	INVX1 INVX1_1689 ( .gnd(gnd), .vdd(vdd), .A(_10218_), .Y(_10261_) );
	AOI22X1 AOI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_msip), .B(_10261_), .C(csr_gpr_iu_csr_mtval_3_), .D(_8618__bF_buf0), .Y(_10262_) );
	OAI21X1 OAI21X1_4244 ( .gnd(gnd), .vdd(vdd), .A(_8864_), .B(_8847__bF_buf6), .C(_10262_), .Y(_10263_) );
	NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp0cfg_3_), .B(_8372__bF_buf1), .Y(_10264_) );
	OAI21X1 OAI21X1_4245 ( .gnd(gnd), .vdd(vdd), .A(_8700_), .B(_10215_), .C(_10264_), .Y(_10265_) );
	NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_10265_), .B(_10263_), .Y(_10266_) );
	NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_10260_), .B(_10266_), .C(_10259_), .Y(_10267_) );
	OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_10267_), .B(_10252_), .Y(csr_3_) );
	NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_4_), .B(_10165_), .Y(_10268_) );
	OAI21X1 OAI21X1_4246 ( .gnd(gnd), .vdd(vdd), .A(_9360_), .B(_8061_), .C(_10268_), .Y(_10269_) );
	AOI21X1 AOI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_16_), .B(_9234__bF_buf3), .C(_10269_), .Y(_10270_) );
	OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_4_), .B(csr_gpr_iu_csr_mideleg_4_), .Y(_10271_) );
	OAI22X1 OAI22X1_777 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(_9019__bF_buf4), .C(_6899_), .D(_10162_), .Y(_10272_) );
	AOI21X1 AOI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_10170_), .B(_10271_), .C(_10272_), .Y(_10273_) );
	AOI22X1 AOI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf0), .B(csr_gpr_iu_csr_pmpaddr2_4_), .C(csr_gpr_iu_csr_mtval_4_), .D(_8618__bF_buf6), .Y(_10274_) );
	NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_10270_), .B(_10274_), .C(_10273_), .Y(_10275_) );
	AOI22X1 AOI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_4_), .B(_8117__bF_buf0), .C(csr_gpr_iu_csr_stval_4_), .D(_7960__bF_buf2), .Y(_10276_) );
	AOI22X1 AOI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp4cfg_4_), .B(_8327__bF_buf1), .C(csr_gpr_iu_csr_pmp0cfg_4_), .D(_8372__bF_buf0), .Y(_10277_) );
	AOI22X1 AOI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_4_), .B(_7435__bF_buf4), .C(csr_gpr_iu_csr_mcause_4_), .D(_10235_), .Y(_10278_) );
	AOI22X1 AOI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf0), .B(csr_gpr_iu_csr_sscratch_4_), .C(csr_gpr_iu_csr_pmpaddr1_4_), .D(_8233__bF_buf3), .Y(_10279_) );
	NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_10279_), .B(_10278_), .Y(_10280_) );
	AOI22X1 AOI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_4_), .B(_8846__bF_buf2), .C(csr_gpr_iu_csr_mscratch_4_), .D(_8417__bF_buf1), .Y(_10281_) );
	NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_4_), .B(_7584__bF_buf2), .Y(_10282_) );
	NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_4_), .B(_8280__bF_buf2), .Y(_10283_) );
	NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_10282_), .B(_10283_), .C(_10281_), .Y(_10284_) );
	NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_10280_), .B(_10284_), .Y(_10285_) );
	NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_10276_), .B(_10277_), .C(_10285_), .Y(_10286_) );
	OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_10286_), .B(_10275_), .Y(csr_4_) );
	AOI22X1 AOI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_5_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_5_), .D(_10208_), .Y(_10287_) );
	AOI22X1 AOI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(_10163_), .B(csr_gpr_iu_csr_mtvec_5_), .C(csr_gpr_iu_csr_mscratch_5_), .D(_8417__bF_buf0), .Y(_10288_) );
	AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_10288_), .B(_10287_), .Y(_10289_) );
	AOI22X1 AOI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_5_), .B(_8165__bF_buf0), .C(csr_gpr_iu_csr_scause_5_), .D(_7435__bF_buf3), .Y(_10290_) );
	OAI21X1 OAI21X1_4247 ( .gnd(gnd), .vdd(vdd), .A(_7653_), .B(_7586__bF_buf3), .C(_10290_), .Y(_10291_) );
	AOI21X1 AOI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_5_), .B(_8062__bF_buf1), .C(_10291_), .Y(_10292_) );
	AOI22X1 AOI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_17_), .B(_9234__bF_buf2), .C(csr_gpr_iu_csr_stval_5_), .D(_10199_), .Y(_10293_) );
	OAI21X1 OAI21X1_4248 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_10196_), .C(_10293_), .Y(_10294_) );
	AOI22X1 AOI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stie), .B(_8469_), .C(csr_gpr_iu_csr_spie), .D(_9144_), .Y(_10295_) );
	NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_5_), .B(_8117__bF_buf6), .Y(_10296_) );
	NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_5_), .B(_7319__bF_buf0), .Y(_10297_) );
	NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_10295_), .B(_10297_), .C(_10296_), .Y(_10298_) );
	NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_10294_), .B(_10298_), .Y(_10299_) );
	AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_10299_), .B(_10292_), .Y(_10300_) );
	NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spie), .B(_9110__bF_buf1), .Y(_10301_) );
	AOI22X1 AOI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp0cfg_5_), .B(_8372__bF_buf6), .C(csr_gpr_iu_csr_pmp4cfg_5_), .D(_8327__bF_buf0), .Y(_10302_) );
	OAI21X1 OAI21X1_4249 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_5_), .B(csr_gpr_iu_csr_mideleg_5_), .C(_8489__bF_buf4), .Y(_10303_) );
	NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .B(_10303_), .C(_10302_), .Y(_10304_) );
	NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_5_), .B(_8233__bF_buf2), .Y(_10305_) );
	AOI22X1 AOI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_5_), .B(_8846__bF_buf1), .C(csr_gpr_iu_csr_mcause_5_), .D(_10214_), .Y(_10306_) );
	OAI22X1 OAI22X1_778 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_10218_), .C(_8630_), .D(_8617_), .Y(_10307_) );
	AOI21X1 AOI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_5_), .B(_8280__bF_buf1), .C(_10307_), .Y(_10308_) );
	NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_10305_), .B(_10306_), .C(_10308_), .Y(_10309_) );
	NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_10304_), .B(_10309_), .Y(_10310_) );
	NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_10289_), .B(_10310_), .C(_10300_), .Y(csr_5_) );
	AOI22X1 AOI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_6_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_6_), .D(_10208_), .Y(_10311_) );
	OAI21X1 OAI21X1_4250 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9019__bF_buf3), .C(_10311_), .Y(_10312_) );
	AOI21X1 AOI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_6_), .B(_8417__bF_buf5), .C(_10312_), .Y(_10313_) );
	AOI22X1 AOI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_6_), .B(_10214_), .C(csr_gpr_iu_csr_mtval_6_), .D(_8618__bF_buf5), .Y(_10314_) );
	OAI21X1 OAI21X1_4251 ( .gnd(gnd), .vdd(vdd), .A(_8882_), .B(_8847__bF_buf5), .C(_10314_), .Y(_10315_) );
	NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_6_), .B(_8165__bF_buf4), .Y(_10316_) );
	OAI21X1 OAI21X1_4252 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_6_), .B(csr_gpr_iu_csr_mideleg_6_), .C(_8489__bF_buf3), .Y(_10317_) );
	NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_10316_), .B(_10317_), .Y(_10318_) );
	NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_10318_), .B(_10315_), .Y(_10319_) );
	AOI22X1 AOI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .B(csr_gpr_iu_csr_sscratch_6_), .C(csr_gpr_iu_csr_sepc_6_), .D(_7584__bF_buf1), .Y(_10320_) );
	AOI22X1 AOI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_6_), .B(_8062__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr3_6_), .D(_8117__bF_buf5), .Y(_10321_) );
	NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_10320_), .B(_10321_), .Y(_10322_) );
	INVX1 INVX1_1690 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_6_), .Y(_10323_) );
	NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_6_), .B(_8233__bF_buf1), .Y(_10324_) );
	OAI21X1 OAI21X1_4253 ( .gnd(gnd), .vdd(vdd), .A(_10323_), .B(_8279_), .C(_10324_), .Y(_10325_) );
	AOI21X1 AOI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp4cfg_6_), .B(_8327__bF_buf6), .C(_10325_), .Y(_10326_) );
	AOI22X1 AOI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf2), .B(csr_gpr_iu_csr_scause_6_), .C(csr_gpr_iu_csr_stval_6_), .D(_10199_), .Y(_10327_) );
	AOI22X1 AOI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf1), .B(biu_mmu_ag0_18_), .C(csr_gpr_iu_csr_pmp0cfg_6_), .D(_8372__bF_buf5), .Y(_10328_) );
	NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(_10327_), .B(_10328_), .C(_10326_), .Y(_10329_) );
	NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_10322_), .B(_10329_), .Y(_10330_) );
	NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .B(_10319_), .C(_10330_), .Y(csr_6_) );
	INVX1 INVX1_1691 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_7_), .Y(_10331_) );
	AOI22X1 AOI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtie), .B(_10244_), .C(csr_gpr_iu_csr_mscratch_7_), .D(_8417__bF_buf4), .Y(_10332_) );
	OAI21X1 OAI21X1_4254 ( .gnd(gnd), .vdd(vdd), .A(_10331_), .B(_9019__bF_buf2), .C(_10332_), .Y(_10333_) );
	AOI21X1 AOI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_7_), .B(_10186_), .C(_10333_), .Y(_10334_) );
	AOI22X1 AOI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_19_), .B(_9234__bF_buf0), .C(csr_gpr_iu_csr_stval_7_), .D(_10199_), .Y(_10335_) );
	OAI21X1 OAI21X1_4255 ( .gnd(gnd), .vdd(vdd), .A(_7672_), .B(_7586__bF_buf2), .C(_10335_), .Y(_10336_) );
	NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_7_), .B(_8062__bF_buf5), .Y(_10337_) );
	AOI22X1 AOI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_7_), .B(_8165__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_7_), .D(_8117__bF_buf4), .Y(_10338_) );
	AOI22X1 AOI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf3), .B(csr_gpr_iu_csr_sscratch_7_), .C(csr_gpr_iu_csr_scause_7_), .D(_7435__bF_buf1), .Y(_10339_) );
	NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_10337_), .B(_10339_), .C(_10338_), .Y(_10340_) );
	NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_10336_), .B(_10340_), .Y(_10341_) );
	OAI22X1 OAI22X1_779 ( .gnd(gnd), .vdd(vdd), .A(_7293_), .B(_10218_), .C(_8634_), .D(_8617_), .Y(_10342_) );
	AOI21X1 AOI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_7_), .B(_10214_), .C(_10342_), .Y(_10343_) );
	OAI21X1 OAI21X1_4256 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_8847__bF_buf4), .C(_10343_), .Y(_10344_) );
	AOI22X1 AOI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_7_), .B(_8233__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr0_7_), .D(_8280__bF_buf0), .Y(_10345_) );
	AOI22X1 AOI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp0cfg_7_), .B(_8372__bF_buf4), .C(csr_gpr_iu_csr_pmp4cfg_7_), .D(_8327__bF_buf5), .Y(_10346_) );
	INVX1 INVX1_1692 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf0), .Y(_10347_) );
	OAI21X1 OAI21X1_4257 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_7_), .B(csr_gpr_iu_csr_mideleg_7_), .C(_8489__bF_buf2), .Y(_10348_) );
	OAI21X1 OAI21X1_4258 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_10347_), .C(_10348_), .Y(_10349_) );
	AOI21X1 AOI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_7_), .B(_10208_), .C(_10349_), .Y(_10350_) );
	NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_10345_), .B(_10346_), .C(_10350_), .Y(_10351_) );
	NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_10344_), .B(_10351_), .Y(_10352_) );
	NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_10334_), .B(_10341_), .C(_10352_), .Y(csr_7_) );
	AOI22X1 AOI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_8_), .B(_7323__bF_buf3), .C(csr_gpr_iu_csr_mtval_8_), .D(_8618__bF_buf4), .Y(_10353_) );
	AOI22X1 AOI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_8_), .B(_7435__bF_buf0), .C(csr_gpr_iu_csr_pmpaddr0_8_), .D(_8280__bF_buf5), .Y(_10354_) );
	NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_10353_), .B(_10354_), .Y(_10355_) );
	NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spp), .B(_9144_), .Y(_10356_) );
	OAI21X1 OAI21X1_4259 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9019__bF_buf1), .C(_10356_), .Y(_10357_) );
	AOI21X1 AOI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_spp), .B(_9110__bF_buf3), .C(_10357_), .Y(_10358_) );
	AOI22X1 AOI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf3), .B(biu_mmu_ag0_20_), .C(csr_gpr_iu_csr_stvec_8_), .D(_8062__bF_buf4), .Y(_10359_) );
	AOI22X1 AOI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(_10227_), .B(csr_gpr_iu_csr_minstret_8_), .C(csr_gpr_iu_csr_mcycle_8_), .D(_10165_), .Y(_10360_) );
	NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_10359_), .B(_10360_), .C(_10358_), .Y(_10361_) );
	NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_10355_), .B(_10361_), .Y(_10362_) );
	AOI22X1 AOI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf0), .B(csr_gpr_iu_csr_sepc_8_), .C(csr_gpr_iu_csr_pmpaddr3_8_), .D(_8117__bF_buf3), .Y(_10363_) );
	OAI21X1 OAI21X1_4260 ( .gnd(gnd), .vdd(vdd), .A(_8890_), .B(_8847__bF_buf3), .C(_10363_), .Y(_10364_) );
	OAI21X1 OAI21X1_4261 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_8_), .B(csr_gpr_iu_csr_mideleg_8_), .C(_10170_), .Y(_10365_) );
	OAI21X1 OAI21X1_4262 ( .gnd(gnd), .vdd(vdd), .A(_7984_), .B(_7959_), .C(_10365_), .Y(_10366_) );
	INVX1 INVX1_1693 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_8_), .Y(_10367_) );
	NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_0_), .B(_8327__bF_buf4), .Y(_10368_) );
	OAI21X1 OAI21X1_4263 ( .gnd(gnd), .vdd(vdd), .A(_10367_), .B(_8232_), .C(_10368_), .Y(_10369_) );
	NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_10369_), .B(_10366_), .Y(_10370_) );
	AOI22X1 AOI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf3), .B(csr_gpr_iu_csr_pmpaddr2_8_), .C(csr_gpr_iu_csr_mcause_8_), .D(_10235_), .Y(_10371_) );
	AOI22X1 AOI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(_8372__bF_buf3), .B(csr_gpr_iu_csr_pmp1cfg_0_), .C(csr_gpr_iu_csr_mscratch_8_), .D(_8417__bF_buf3), .Y(_10372_) );
	NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(_10371_), .B(_10372_), .C(_10370_), .Y(_10373_) );
	NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_10364_), .B(_10373_), .Y(_10374_) );
	NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_10362_), .B(_10374_), .Y(csr_8_) );
	AOI22X1 AOI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seie), .B(_10244_), .C(csr_gpr_iu_csr_minstret_9_), .D(_10208_), .Y(_10375_) );
	OAI21X1 OAI21X1_4264 ( .gnd(gnd), .vdd(vdd), .A(_9538_), .B(_9019__bF_buf0), .C(_10375_), .Y(_10376_) );
	INVX1 INVX1_1694 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_9_), .Y(_10377_) );
	OAI21X1 OAI21X1_4265 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_9_), .B(csr_gpr_iu_csr_mideleg_9_), .C(_8489__bF_buf1), .Y(_10378_) );
	OAI21X1 OAI21X1_4266 ( .gnd(gnd), .vdd(vdd), .A(_10377_), .B(_8116_), .C(_10378_), .Y(_10379_) );
	NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_10379_), .B(_10376_), .Y(_10380_) );
	NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_21_), .B(_9234__bF_buf2), .Y(_10381_) );
	OAI21X1 OAI21X1_4267 ( .gnd(gnd), .vdd(vdd), .A(_7987_), .B(_10198_), .C(_10381_), .Y(_10382_) );
	OAI22X1 OAI22X1_780 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_8061_), .C(_7296_), .D(_10196_), .Y(_10383_) );
	NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_10383_), .B(_10382_), .Y(_10384_) );
	AOI22X1 AOI22X1_506 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_1_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_9_), .D(_8280__bF_buf4), .Y(_10385_) );
	AOI22X1 AOI22X1_507 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seip), .B(_10261_), .C(csr_gpr_iu_csr_pmp1cfg_1_), .D(_8372__bF_buf2), .Y(_10386_) );
	AOI22X1 AOI22X1_508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_9_), .B(_10214_), .C(csr_gpr_iu_csr_mtval_9_), .D(_8618__bF_buf3), .Y(_10387_) );
	OAI21X1 OAI21X1_4268 ( .gnd(gnd), .vdd(vdd), .A(_8897_), .B(_8847__bF_buf2), .C(_10387_), .Y(_10388_) );
	AOI21X1 AOI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_9_), .B(_8417__bF_buf2), .C(_10388_), .Y(_10389_) );
	NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_10385_), .B(_10386_), .C(_10389_), .Y(_10390_) );
	AOI22X1 AOI22X1_509 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf6), .B(csr_gpr_iu_csr_scause_9_), .C(csr_gpr_iu_csr_pmpaddr1_9_), .D(_8233__bF_buf5), .Y(_10391_) );
	OAI21X1 OAI21X1_4269 ( .gnd(gnd), .vdd(vdd), .A(_7697_), .B(_7586__bF_buf1), .C(_10391_), .Y(_10392_) );
	AOI21X1 AOI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_9_), .B(_7319__bF_buf2), .C(_10392_), .Y(_10393_) );
	NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_9_), .B(_8165__bF_buf2), .Y(_10394_) );
	NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(_7309__bF_buf0), .Y(_10395_) );
	AOI22X1 AOI22X1_510 ( .gnd(gnd), .vdd(vdd), .A(_10186_), .B(csr_gpr_iu_csr_mcycle_9_), .C(csr_gpr_iu_csr_seie), .D(_10395_), .Y(_10396_) );
	NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_10394_), .B(_10396_), .C(_10393_), .Y(_10397_) );
	NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_10397_), .B(_10390_), .Y(_10398_) );
	NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_10380_), .B(_10384_), .C(_10398_), .Y(csr_9_) );
	OAI22X1 OAI22X1_781 ( .gnd(gnd), .vdd(vdd), .A(_9545_), .B(_9019__bF_buf5), .C(_6812_), .D(_10164_), .Y(_10399_) );
	AOI21X1 AOI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_10_), .B(_10227_), .C(_10399_), .Y(_10400_) );
	AOI22X1 AOI22X1_511 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf1), .B(biu_mmu_ag0_22_), .C(csr_gpr_iu_csr_stvec_10_), .D(_8062__bF_buf3), .Y(_10401_) );
	OAI21X1 OAI21X1_4270 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8684__bF_buf1), .C(_10401_), .Y(_10402_) );
	INVX1 INVX1_1695 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_10_), .Y(_10403_) );
	OAI21X1 OAI21X1_4271 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_10_), .B(csr_gpr_iu_csr_mideleg_10_), .C(_10170_), .Y(_10404_) );
	OAI21X1 OAI21X1_4272 ( .gnd(gnd), .vdd(vdd), .A(_10403_), .B(_8279_), .C(_10404_), .Y(_10405_) );
	NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10405_), .Y(_10406_) );
	AOI22X1 AOI22X1_512 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf1), .B(csr_gpr_iu_csr_sscratch_10_), .C(csr_gpr_iu_csr_sepc_10_), .D(_7584__bF_buf5), .Y(_10407_) );
	AOI22X1 AOI22X1_513 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_2_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_mscratch_10_), .D(_8417__bF_buf1), .Y(_10408_) );
	NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_10407_), .B(_10408_), .Y(_10409_) );
	NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_10_), .B(_8233__bF_buf4), .Y(_10410_) );
	OAI21X1 OAI21X1_4273 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8617_), .C(_10410_), .Y(_10411_) );
	OAI22X1 OAI22X1_782 ( .gnd(gnd), .vdd(vdd), .A(_8902_), .B(_8847__bF_buf1), .C(_7476_), .D(_7437_), .Y(_10412_) );
	NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_10412_), .B(_10411_), .Y(_10413_) );
	AOI22X1 AOI22X1_514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_10_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_stval_10_), .D(_7960__bF_buf1), .Y(_10414_) );
	AOI22X1 AOI22X1_515 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr2_10_), .C(csr_gpr_iu_csr_pmp1cfg_2_), .D(_8372__bF_buf1), .Y(_10415_) );
	NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_10414_), .B(_10415_), .C(_10413_), .Y(_10416_) );
	NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .B(_10416_), .Y(_10417_) );
	NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_10400_), .B(_10406_), .C(_10417_), .Y(csr_10_) );
	AOI22X1 AOI22X1_516 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meie), .B(_10244_), .C(csr_gpr_iu_csr_mscratch_11_), .D(_8417__bF_buf0), .Y(_10418_) );
	OAI21X1 OAI21X1_4274 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_9019__bF_buf4), .C(_10418_), .Y(_10419_) );
	AOI21X1 AOI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_11_), .B(_10186_), .C(_10419_), .Y(_10420_) );
	AOI22X1 AOI22X1_517 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_23_), .B(_9234__bF_buf0), .C(csr_gpr_iu_csr_stval_11_), .D(_10199_), .Y(_10421_) );
	AOI22X1 AOI22X1_518 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf4), .B(csr_gpr_iu_csr_sepc_11_), .C(csr_gpr_iu_csr_scause_11_), .D(_7435__bF_buf5), .Y(_10422_) );
	NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_10422_), .B(_10421_), .Y(_10423_) );
	AOI22X1 AOI22X1_519 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_11_), .B(_7319__bF_buf0), .C(csr_gpr_iu_csr_stvec_11_), .D(_8062__bF_buf2), .Y(_10424_) );
	AOI22X1 AOI22X1_520 ( .gnd(gnd), .vdd(vdd), .A(_8117__bF_buf1), .B(csr_gpr_iu_csr_pmpaddr3_11_), .C(csr_gpr_iu_csr_pmpaddr2_11_), .D(_10182__bF_buf1), .Y(_10425_) );
	NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10425_), .Y(_10426_) );
	NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_10423_), .B(_10426_), .Y(_10427_) );
	AOI22X1 AOI22X1_521 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip), .B(_10261_), .C(csr_gpr_iu_csr_mtval_11_), .D(_8618__bF_buf2), .Y(_10428_) );
	OAI21X1 OAI21X1_4275 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8847__bF_buf0), .C(_10428_), .Y(_10429_) );
	AOI21X1 AOI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_11_), .B(_10214_), .C(_10429_), .Y(_10430_) );
	NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_3_), .B(_8327__bF_buf1), .Y(_10431_) );
	NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp1cfg_3_), .B(_8372__bF_buf0), .Y(_10432_) );
	AOI22X1 AOI22X1_522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_11_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_11_), .D(_8280__bF_buf3), .Y(_10433_) );
	NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .B(_10432_), .C(_10433_), .Y(_10434_) );
	NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_0_), .B(_9110__bF_buf2), .Y(_10435_) );
	OAI21X1 OAI21X1_4276 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_11_), .B(csr_gpr_iu_csr_mideleg_11_), .C(_8489__bF_buf0), .Y(_10436_) );
	AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10435_), .Y(_10437_) );
	OAI21X1 OAI21X1_4277 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(_10209_), .C(_10437_), .Y(_10438_) );
	NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_10438_), .B(_10434_), .Y(_10439_) );
	AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_10439_), .B(_10430_), .Y(_10440_) );
	NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10427_), .C(_10440_), .Y(csr_11_) );
	NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_12_), .B(_8618__bF_buf1), .Y(_10441_) );
	AOI22X1 AOI22X1_523 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf3), .B(csr_gpr_iu_csr_sepc_12_), .C(csr_gpr_iu_csr_scause_12_), .D(_7435__bF_buf4), .Y(_10442_) );
	AOI22X1 AOI22X1_524 ( .gnd(gnd), .vdd(vdd), .A(_10214_), .B(csr_gpr_iu_csr_mcause_12_), .C(csr_gpr_iu_csr_pmpaddr0_12_), .D(_8280__bF_buf2), .Y(_10443_) );
	NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_10442_), .B(_10441_), .C(_10443_), .Y(_10444_) );
	NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_12_), .B(_10163_), .Y(_10445_) );
	NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mpp_1_), .B(_9110__bF_buf1), .Y(_10446_) );
	AOI22X1 AOI22X1_525 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_12_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_12_), .D(_10208_), .Y(_10447_) );
	NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_10445_), .B(_10446_), .C(_10447_), .Y(_10448_) );
	NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_10448_), .B(_10444_), .Y(_10449_) );
	AOI22X1 AOI22X1_526 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_12_), .B(_8165__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_12_), .D(_8117__bF_buf0), .Y(_10450_) );
	OAI21X1 OAI21X1_4278 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_9161__bF_buf3), .C(_10450_), .Y(_10451_) );
	AOI22X1 AOI22X1_527 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_12_), .B(_8062__bF_buf1), .C(csr_gpr_iu_csr_sscratch_12_), .D(_7319__bF_buf4), .Y(_10452_) );
	OAI21X1 OAI21X1_4279 ( .gnd(gnd), .vdd(vdd), .A(_7996_), .B(_10198_), .C(_10452_), .Y(_10453_) );
	NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_10453_), .B(_10451_), .Y(_10454_) );
	AOI22X1 AOI22X1_528 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_4_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_pmp1cfg_4_), .D(_8372__bF_buf6), .Y(_10455_) );
	OAI21X1 OAI21X1_4280 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_12_), .B(csr_gpr_iu_csr_mideleg_12_), .C(_8489__bF_buf5), .Y(_10456_) );
	NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_10456_), .B(_10455_), .Y(_10457_) );
	INVX1 INVX1_1696 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_12_), .Y(_10458_) );
	AOI22X1 AOI22X1_529 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_12_), .B(_8846__bF_buf0), .C(csr_gpr_iu_csr_mscratch_12_), .D(_8417__bF_buf5), .Y(_10459_) );
	OAI21X1 OAI21X1_4281 ( .gnd(gnd), .vdd(vdd), .A(_10458_), .B(_8232_), .C(_10459_), .Y(_10460_) );
	NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_10457_), .B(_10460_), .Y(_10461_) );
	NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_10454_), .B(_10461_), .C(_10449_), .Y(csr_12_) );
	AOI22X1 AOI22X1_530 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_13_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_13_), .D(_10208_), .Y(_10462_) );
	OAI21X1 OAI21X1_4282 ( .gnd(gnd), .vdd(vdd), .A(_9049_), .B(_9019__bF_buf3), .C(_10462_), .Y(_10463_) );
	AOI21X1 AOI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_13_), .B(_8417__bF_buf4), .C(_10463_), .Y(_10464_) );
	AOI22X1 AOI22X1_531 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_13_), .B(_10214_), .C(csr_gpr_iu_csr_mtval_13_), .D(_8618__bF_buf0), .Y(_10465_) );
	OAI21X1 OAI21X1_4283 ( .gnd(gnd), .vdd(vdd), .A(_8918_), .B(_8847__bF_buf7), .C(_10465_), .Y(_10466_) );
	OAI21X1 OAI21X1_4284 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_13_), .B(csr_gpr_iu_csr_mideleg_13_), .C(_8489__bF_buf4), .Y(_10467_) );
	OAI21X1 OAI21X1_4285 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_8162__bF_buf1), .C(_10467_), .Y(_10468_) );
	NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_10468_), .B(_10466_), .Y(_10469_) );
	NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_10464_), .B(_10469_), .Y(_10470_) );
	AOI22X1 AOI22X1_532 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf3), .B(csr_gpr_iu_csr_sscratch_13_), .C(csr_gpr_iu_csr_sepc_13_), .D(_7584__bF_buf2), .Y(_10471_) );
	OAI21X1 OAI21X1_4286 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .B(_8061_), .C(_10471_), .Y(_10472_) );
	OAI22X1 OAI22X1_783 ( .gnd(gnd), .vdd(vdd), .A(_8403_), .B(_8371_), .C(_8132_), .D(_8116_), .Y(_10473_) );
	NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_10473_), .B(_10472_), .Y(_10474_) );
	OAI22X1 OAI22X1_784 ( .gnd(gnd), .vdd(vdd), .A(_7488_), .B(_7437_), .C(_7999_), .D(_10198_), .Y(_10475_) );
	AOI21X1 AOI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_ag0_25_), .B(_9234__bF_buf3), .C(_10475_), .Y(_10476_) );
	OAI22X1 OAI22X1_785 ( .gnd(gnd), .vdd(vdd), .A(_8295_), .B(_8279_), .C(_8249_), .D(_8232_), .Y(_10477_) );
	AOI21X1 AOI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_5_), .B(_8327__bF_buf6), .C(_10477_), .Y(_10478_) );
	NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10476_), .C(_10474_), .Y(_10479_) );
	OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_10470_), .B(_10479_), .Y(csr_13_) );
	AOI22X1 AOI22X1_533 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_14_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_14_), .D(_10208_), .Y(_10480_) );
	OAI21X1 OAI21X1_4287 ( .gnd(gnd), .vdd(vdd), .A(_9669_), .B(_9019__bF_buf2), .C(_10480_), .Y(_10481_) );
	AOI21X1 AOI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_14_), .B(_8417__bF_buf3), .C(_10481_), .Y(_10482_) );
	AOI22X1 AOI22X1_534 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_14_), .B(_10214_), .C(csr_gpr_iu_csr_mtval_14_), .D(_8618__bF_buf6), .Y(_10483_) );
	OAI21X1 OAI21X1_4288 ( .gnd(gnd), .vdd(vdd), .A(_8927_), .B(_8847__bF_buf6), .C(_10483_), .Y(_10484_) );
	INVX1 INVX1_1697 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_14_), .Y(_10485_) );
	OAI21X1 OAI21X1_4289 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_14_), .B(csr_gpr_iu_csr_mideleg_14_), .C(_8489__bF_buf3), .Y(_10486_) );
	OAI21X1 OAI21X1_4290 ( .gnd(gnd), .vdd(vdd), .A(_10485_), .B(_8162__bF_buf0), .C(_10486_), .Y(_10487_) );
	NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_10487_), .B(_10484_), .Y(_10488_) );
	NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_10482_), .B(_10488_), .Y(_10489_) );
	AOI22X1 AOI22X1_535 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf2), .B(csr_gpr_iu_csr_sscratch_14_), .C(csr_gpr_iu_csr_sepc_14_), .D(_7584__bF_buf1), .Y(_10490_) );
	OAI21X1 OAI21X1_4291 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_8061_), .C(_10490_), .Y(_10491_) );
	AOI21X1 AOI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_14_), .B(_8117__bF_buf6), .C(_10491_), .Y(_10492_) );
	INVX1 INVX1_1698 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_14_), .Y(_10493_) );
	NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_14_), .B(_8233__bF_buf2), .Y(_10494_) );
	OAI21X1 OAI21X1_4292 ( .gnd(gnd), .vdd(vdd), .A(_10493_), .B(_8279_), .C(_10494_), .Y(_10495_) );
	AOI21X1 AOI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_6_), .B(_8327__bF_buf5), .C(_10495_), .Y(_10496_) );
	AOI22X1 AOI22X1_536 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf3), .B(csr_gpr_iu_csr_scause_14_), .C(csr_gpr_iu_csr_stval_14_), .D(_10199_), .Y(_10497_) );
	AOI22X1 AOI22X1_537 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf2), .B(biu_mmu_ag0_26_), .C(csr_gpr_iu_csr_pmp1cfg_6_), .D(_8372__bF_buf5), .Y(_10498_) );
	AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_10498_), .B(_10497_), .Y(_10499_) );
	NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(_10492_), .B(_10499_), .C(_10496_), .Y(_10500_) );
	OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_10489_), .B(_10500_), .Y(csr_14_) );
	NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_15_), .B(_10186_), .Y(_10501_) );
	OAI21X1 OAI21X1_4293 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_10209_), .C(_10501_), .Y(_10502_) );
	AOI21X1 AOI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_15_), .B(_10163_), .C(_10502_), .Y(_10503_) );
	OAI21X1 OAI21X1_4294 ( .gnd(gnd), .vdd(vdd), .A(_8436_), .B(_8416_), .C(_10503_), .Y(_10504_) );
	OAI22X1 OAI22X1_786 ( .gnd(gnd), .vdd(vdd), .A(_8650_), .B(_8617_), .C(_8760_), .D(_10215_), .Y(_10505_) );
	AOI21X1 AOI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_15_), .B(_8846__bF_buf3), .C(_10505_), .Y(_10506_) );
	NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_15_), .B(_8165__bF_buf0), .Y(_10507_) );
	OAI21X1 OAI21X1_4295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_15_), .B(csr_gpr_iu_csr_mideleg_15_), .C(_8489__bF_buf2), .Y(_10508_) );
	NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(_10507_), .B(_10508_), .C(_10506_), .Y(_10509_) );
	NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_10504_), .B(_10509_), .Y(_10510_) );
	OAI22X1 OAI22X1_787 ( .gnd(gnd), .vdd(vdd), .A(_7372_), .B(_7320__bF_buf1), .C(_7765_), .D(_7586__bF_buf0), .Y(_10511_) );
	AOI21X1 AOI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_15_), .B(_8117__bF_buf5), .C(_10511_), .Y(_10512_) );
	OAI21X1 OAI21X1_4296 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_8061_), .C(_10512_), .Y(_10513_) );
	OAI22X1 OAI22X1_788 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8279_), .C(_8252_), .D(_8232_), .Y(_10514_) );
	AOI21X1 AOI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp5cfg_7_), .B(_8327__bF_buf4), .C(_10514_), .Y(_10515_) );
	AOI22X1 AOI22X1_538 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf2), .B(csr_gpr_iu_csr_scause_15_), .C(csr_gpr_iu_csr_stval_15_), .D(_10199_), .Y(_10516_) );
	AOI22X1 AOI22X1_539 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf1), .B(biu_mmu_ag0_27_), .C(csr_gpr_iu_csr_pmp1cfg_7_), .D(_8372__bF_buf4), .Y(_10517_) );
	NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_10516_), .B(_10517_), .C(_10515_), .Y(_10518_) );
	NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_10518_), .B(_10513_), .Y(_10519_) );
	NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_10510_), .B(_10519_), .Y(csr_15_) );
	OAI22X1 OAI22X1_789 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9019__bF_buf1), .C(_7185_), .D(_10164_), .Y(_10520_) );
	AOI21X1 AOI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_16_), .B(_10227_), .C(_10520_), .Y(_10521_) );
	AOI22X1 AOI22X1_540 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf0), .B(biu_mmu_ag0_28_), .C(csr_gpr_iu_csr_stvec_16_), .D(_8062__bF_buf0), .Y(_10522_) );
	OAI21X1 OAI21X1_4297 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_8684__bF_buf0), .C(_10522_), .Y(_10523_) );
	OAI21X1 OAI21X1_4298 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_16_), .B(csr_gpr_iu_csr_mideleg_16_), .C(_10170_), .Y(_10524_) );
	OAI21X1 OAI21X1_4299 ( .gnd(gnd), .vdd(vdd), .A(_8008_), .B(_7959_), .C(_10524_), .Y(_10525_) );
	NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_10523_), .B(_10525_), .Y(_10526_) );
	AOI22X1 AOI22X1_541 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf1), .B(csr_gpr_iu_csr_sscratch_16_), .C(csr_gpr_iu_csr_sepc_16_), .D(_7584__bF_buf0), .Y(_10527_) );
	NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_16_), .B(_8280__bF_buf1), .Y(_10528_) );
	NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_16_), .B(_8417__bF_buf2), .Y(_10529_) );
	NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_10527_), .B(_10529_), .C(_10528_), .Y(_10530_) );
	AOI22X1 AOI22X1_542 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_16_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_mtval_16_), .D(_8618__bF_buf5), .Y(_10531_) );
	AOI22X1 AOI22X1_543 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_16_), .B(_8846__bF_buf2), .C(csr_gpr_iu_csr_pmp2cfg_0_), .D(_8372__bF_buf3), .Y(_10532_) );
	AOI22X1 AOI22X1_544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_16_), .B(_7435__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_16_), .D(_8117__bF_buf4), .Y(_10533_) );
	AOI22X1 AOI22X1_545 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_0_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_16_), .D(_10182__bF_buf0), .Y(_10534_) );
	AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_10533_), .B(_10534_), .Y(_10535_) );
	NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(_10531_), .B(_10532_), .C(_10535_), .Y(_10536_) );
	NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_10530_), .B(_10536_), .Y(_10537_) );
	NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(_10521_), .B(_10526_), .C(_10537_), .Y(csr_16_) );
	AOI22X1 AOI22X1_546 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf5), .B(csr_gpr_iu_csr_sepc_17_), .C(csr_gpr_iu_csr_scause_17_), .D(_7435__bF_buf0), .Y(_10538_) );
	OAI21X1 OAI21X1_4300 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_8617_), .C(_10538_), .Y(_10539_) );
	OAI22X1 OAI22X1_790 ( .gnd(gnd), .vdd(vdd), .A(_8301_), .B(_8279_), .C(_8770_), .D(_10215_), .Y(_10540_) );
	NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_10540_), .B(_10539_), .Y(_10541_) );
	AOI22X1 AOI22X1_547 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf0), .B(csr_gpr_iu_csr_mprv), .C(csr_gpr_iu_csr_mcycle_17_), .D(_10186_), .Y(_10542_) );
	OAI21X1 OAI21X1_4301 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_9019__bF_buf0), .C(_10542_), .Y(_10543_) );
	AOI21X1 AOI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_17_), .B(_10208_), .C(_10543_), .Y(_10544_) );
	AOI22X1 AOI22X1_548 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_17_), .B(_8165__bF_buf4), .C(csr_gpr_iu_csr_pmpaddr3_17_), .D(_8117__bF_buf3), .Y(_10545_) );
	OAI21X1 OAI21X1_4302 ( .gnd(gnd), .vdd(vdd), .A(_9199_), .B(_9161__bF_buf2), .C(_10545_), .Y(_10546_) );
	AOI22X1 AOI22X1_549 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_17_), .B(_7319__bF_buf0), .C(csr_gpr_iu_csr_stval_17_), .D(_10199_), .Y(_10547_) );
	OAI21X1 OAI21X1_4303 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_8061_), .C(_10547_), .Y(_10548_) );
	OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_10546_), .B(_10548_), .Y(_10549_) );
	AOI22X1 AOI22X1_550 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_1_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmp2cfg_1_), .D(_8372__bF_buf2), .Y(_10550_) );
	OAI21X1 OAI21X1_4304 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_17_), .B(csr_gpr_iu_csr_mideleg_17_), .C(_8489__bF_buf1), .Y(_10551_) );
	OAI22X1 OAI22X1_791 ( .gnd(gnd), .vdd(vdd), .A(_8440_), .B(_8416_), .C(_8941_), .D(_8847__bF_buf5), .Y(_10552_) );
	AOI21X1 AOI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_17_), .B(_8233__bF_buf0), .C(_10552_), .Y(_10553_) );
	NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(_10550_), .B(_10551_), .C(_10553_), .Y(_10554_) );
	NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_10554_), .B(_10549_), .Y(_10555_) );
	NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(_10541_), .B(_10544_), .C(_10555_), .Y(csr_17_) );
	AOI22X1 AOI22X1_551 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .B(csr_gpr_iu_csr_sscratch_18_), .C(csr_gpr_iu_csr_sepc_18_), .D(_7584__bF_buf4), .Y(_10556_) );
	AOI22X1 AOI22X1_552 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf3), .B(csr_gpr_iu_csr_pmpaddr2_18_), .C(csr_gpr_iu_csr_mcause_18_), .D(_10235_), .Y(_10557_) );
	AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_10557_), .B(_10556_), .Y(_10558_) );
	AOI22X1 AOI22X1_553 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_sum), .B(_9110__bF_buf3), .C(biu_mmu_ag0_30_), .D(_9234__bF_buf3), .Y(_10559_) );
	OAI21X1 OAI21X1_4305 ( .gnd(gnd), .vdd(vdd), .A(_6996_), .B(_10162_), .C(_10559_), .Y(_10560_) );
	AOI22X1 AOI22X1_554 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_18_), .B(_8062__bF_buf5), .C(biu_mmu_sum), .D(_9144_), .Y(_10561_) );
	AOI22X1 AOI22X1_555 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_18_), .B(_10163_), .C(csr_gpr_iu_csr_mcycle_18_), .D(_10165_), .Y(_10562_) );
	NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_10561_), .B(_10562_), .Y(_10563_) );
	NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_10560_), .B(_10563_), .Y(_10564_) );
	AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_10564_), .B(_10558_), .Y(_10565_) );
	NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp2cfg_2_), .B(_8372__bF_buf1), .Y(_10566_) );
	OAI21X1 OAI21X1_4306 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_7437_), .C(_10566_), .Y(_10567_) );
	AOI21X1 AOI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_18_), .B(_8846__bF_buf1), .C(_10567_), .Y(_10568_) );
	AOI22X1 AOI22X1_556 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtval_18_), .B(_8618__bF_buf4), .C(csr_gpr_iu_csr_stval_18_), .D(_7960__bF_buf0), .Y(_10569_) );
	NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_18_), .B(_8417__bF_buf1), .Y(_10570_) );
	OAI21X1 OAI21X1_4307 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_18_), .B(csr_gpr_iu_csr_mideleg_18_), .C(_10170_), .Y(_10571_) );
	NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_10570_), .B(_10571_), .C(_10569_), .Y(_10572_) );
	NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_2_), .B(_8327__bF_buf1), .Y(_10573_) );
	NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_18_), .B(_8233__bF_buf5), .Y(_10574_) );
	AOI22X1 AOI22X1_557 ( .gnd(gnd), .vdd(vdd), .A(_8117__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr3_18_), .C(csr_gpr_iu_csr_pmpaddr0_18_), .D(_8280__bF_buf0), .Y(_10575_) );
	NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_10573_), .B(_10574_), .C(_10575_), .Y(_10576_) );
	NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_10576_), .B(_10572_), .Y(_10577_) );
	NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_10568_), .B(_10577_), .C(_10565_), .Y(csr_18_) );
	OAI22X1 OAI22X1_792 ( .gnd(gnd), .vdd(vdd), .A(_7808_), .B(_7586__bF_buf5), .C(_7384_), .D(_9233_), .Y(_10578_) );
	OAI22X1 OAI22X1_793 ( .gnd(gnd), .vdd(vdd), .A(_8390_), .B(_8371_), .C(_8658_), .D(_8617_), .Y(_10579_) );
	NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_10579_), .B(_10578_), .Y(_10580_) );
	OAI22X1 OAI22X1_794 ( .gnd(gnd), .vdd(vdd), .A(_8086_), .B(_8061_), .C(_9147_), .D(_10347_), .Y(_10581_) );
	AOI21X1 AOI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_10227_), .B(csr_gpr_iu_csr_minstret_19_), .C(_10581_), .Y(_10582_) );
	OAI22X1 OAI22X1_795 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_9161__bF_buf1), .C(_6790_), .D(_10164_), .Y(_10583_) );
	NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_mxr), .B(_9144_), .Y(_10584_) );
	OAI21X1 OAI21X1_4308 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_9019__bF_buf5), .C(_10584_), .Y(_10585_) );
	NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_10583_), .B(_10585_), .Y(_10586_) );
	AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_10586_), .B(_10582_), .Y(_10587_) );
	AOI22X1 AOI22X1_558 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf6), .B(csr_gpr_iu_csr_scause_19_), .C(csr_gpr_iu_csr_stval_19_), .D(_10199_), .Y(_10588_) );
	OAI21X1 OAI21X1_4309 ( .gnd(gnd), .vdd(vdd), .A(_8258_), .B(_8232_), .C(_10588_), .Y(_10589_) );
	OAI22X1 OAI22X1_796 ( .gnd(gnd), .vdd(vdd), .A(_8304_), .B(_8279_), .C(_8952_), .D(_8847__bF_buf4), .Y(_10590_) );
	OAI21X1 OAI21X1_4310 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_19_), .B(csr_gpr_iu_csr_mideleg_19_), .C(_10170_), .Y(_10591_) );
	OAI21X1 OAI21X1_4311 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .B(_8116_), .C(_10591_), .Y(_10592_) );
	NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_10590_), .B(_10592_), .Y(_10593_) );
	AOI22X1 AOI22X1_559 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr2_19_), .C(csr_gpr_iu_csr_mscratch_19_), .D(_8417__bF_buf0), .Y(_10594_) );
	AOI22X1 AOI22X1_560 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_3_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_mcause_19_), .D(_10235_), .Y(_10595_) );
	NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_10594_), .B(_10595_), .C(_10593_), .Y(_10596_) );
	NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_10589_), .B(_10596_), .Y(_10597_) );
	NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(_10580_), .B(_10587_), .C(_10597_), .Y(csr_19_) );
	OAI22X1 OAI22X1_797 ( .gnd(gnd), .vdd(vdd), .A(_7819_), .B(_7586__bF_buf4), .C(_7521_), .D(_7437_), .Y(_10598_) );
	AOI21X1 AOI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_20_), .B(_10214_), .C(_10598_), .Y(_10599_) );
	AOI22X1 AOI22X1_561 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_20_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_mtval_20_), .D(_8618__bF_buf3), .Y(_10600_) );
	NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_10600_), .B(_10599_), .Y(_10601_) );
	NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_20_), .B(_10163_), .Y(_10602_) );
	AOI22X1 AOI22X1_562 ( .gnd(gnd), .vdd(vdd), .A(_9110__bF_buf2), .B(csr_gpr_iu_csr_tvm), .C(csr_gpr_iu_csr_mcycle_20_), .D(_10186_), .Y(_10603_) );
	AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_10603_), .B(_10602_), .Y(_10604_) );
	OAI21X1 OAI21X1_4312 ( .gnd(gnd), .vdd(vdd), .A(_7004_), .B(_10209_), .C(_10604_), .Y(_10605_) );
	NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_10605_), .B(_10601_), .Y(_10606_) );
	AOI22X1 AOI22X1_563 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_20_), .B(_8165__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_20_), .D(_8117__bF_buf1), .Y(_10607_) );
	OAI21X1 OAI21X1_4313 ( .gnd(gnd), .vdd(vdd), .A(_9205_), .B(_9161__bF_buf0), .C(_10607_), .Y(_10608_) );
	AOI22X1 AOI22X1_564 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_20_), .B(_8062__bF_buf4), .C(csr_gpr_iu_csr_sscratch_20_), .D(_7319__bF_buf3), .Y(_10609_) );
	OAI21X1 OAI21X1_4314 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_10198_), .C(_10609_), .Y(_10610_) );
	OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_10608_), .B(_10610_), .Y(_10611_) );
	AOI22X1 AOI22X1_565 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_4_), .B(_8327__bF_buf6), .C(csr_gpr_iu_csr_pmp2cfg_4_), .D(_8372__bF_buf0), .Y(_10612_) );
	OAI21X1 OAI21X1_4315 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_20_), .B(csr_gpr_iu_csr_mideleg_20_), .C(_8489__bF_buf0), .Y(_10613_) );
	NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_20_), .B(_8417__bF_buf5), .Y(_10614_) );
	OAI21X1 OAI21X1_4316 ( .gnd(gnd), .vdd(vdd), .A(_8957_), .B(_8847__bF_buf3), .C(_10614_), .Y(_10615_) );
	AOI21X1 AOI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_20_), .B(_8280__bF_buf5), .C(_10615_), .Y(_10616_) );
	NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(_10612_), .B(_10613_), .C(_10616_), .Y(_10617_) );
	NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_10611_), .B(_10617_), .Y(_10618_) );
	NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_10606_), .B(_10618_), .Y(csr_20_) );
	AOI22X1 AOI22X1_566 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_21_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_21_), .D(_10208_), .Y(_10619_) );
	OAI21X1 OAI21X1_4317 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9019__bF_buf4), .C(_10619_), .Y(_10620_) );
	AOI21X1 AOI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_21_), .B(_8417__bF_buf4), .C(_10620_), .Y(_10621_) );
	OAI22X1 OAI22X1_798 ( .gnd(gnd), .vdd(vdd), .A(_8662_), .B(_8617_), .C(_8790_), .D(_10215_), .Y(_10622_) );
	AOI21X1 AOI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_21_), .B(_8846__bF_buf0), .C(_10622_), .Y(_10623_) );
	NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_8532_), .B(_8590_), .Y(_10624_) );
	AOI22X1 AOI22X1_567 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr2_21_), .C(_8489__bF_buf5), .D(_10624_), .Y(_10625_) );
	NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(_10625_), .B(_10623_), .C(_10621_), .Y(_10626_) );
	AOI22X1 AOI22X1_568 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf2), .B(csr_gpr_iu_csr_sscratch_21_), .C(csr_gpr_iu_csr_sepc_21_), .D(_7584__bF_buf3), .Y(_10627_) );
	OAI21X1 OAI21X1_4318 ( .gnd(gnd), .vdd(vdd), .A(_8144_), .B(_8116_), .C(_10627_), .Y(_10628_) );
	AOI21X1 AOI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_21_), .B(_8062__bF_buf3), .C(_10628_), .Y(_10629_) );
	OAI22X1 OAI22X1_799 ( .gnd(gnd), .vdd(vdd), .A(_8307_), .B(_8279_), .C(_8261_), .D(_8232_), .Y(_10630_) );
	AOI21X1 AOI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_5_), .B(_8327__bF_buf5), .C(_10630_), .Y(_10631_) );
	OAI22X1 OAI22X1_800 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_10198_), .C(_7525_), .D(_7437_), .Y(_10632_) );
	OAI22X1 OAI22X1_801 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_9161__bF_buf4), .C(_8393_), .D(_8371_), .Y(_10633_) );
	NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_10632_), .Y(_10634_) );
	NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10634_), .C(_10629_), .Y(_10635_) );
	OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_10635_), .B(_10626_), .Y(csr_21_) );
	AOI22X1 AOI22X1_569 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp6cfg_6_), .B(_8327__bF_buf4), .C(csr_gpr_iu_csr_pmp2cfg_6_), .D(_8372__bF_buf6), .Y(_10636_) );
	OAI21X1 OAI21X1_4319 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_22_), .B(csr_gpr_iu_csr_mideleg_22_), .C(_8489__bF_buf4), .Y(_10637_) );
	NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_10637_), .B(_10636_), .Y(_10638_) );
	INVX1 INVX1_1699 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_tsr), .Y(_10639_) );
	NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_22_), .B(_10186_), .Y(_10640_) );
	OAI21X1 OAI21X1_4320 ( .gnd(gnd), .vdd(vdd), .A(_10639_), .B(_10347_), .C(_10640_), .Y(_10641_) );
	AOI21X1 AOI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_22_), .B(_10163_), .C(_10641_), .Y(_10642_) );
	OAI21X1 OAI21X1_4321 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_10209_), .C(_10642_), .Y(_10643_) );
	NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_10638_), .B(_10643_), .Y(_10644_) );
	AOI22X1 AOI22X1_570 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr2_22_), .B(_8165__bF_buf1), .C(csr_gpr_iu_csr_pmpaddr3_22_), .D(_8117__bF_buf0), .Y(_10645_) );
	OAI21X1 OAI21X1_4322 ( .gnd(gnd), .vdd(vdd), .A(_9210_), .B(_9161__bF_buf3), .C(_10645_), .Y(_10646_) );
	AOI22X1 AOI22X1_571 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_22_), .B(_8062__bF_buf2), .C(csr_gpr_iu_csr_sscratch_22_), .D(_7319__bF_buf1), .Y(_10647_) );
	OAI21X1 OAI21X1_4323 ( .gnd(gnd), .vdd(vdd), .A(_8026_), .B(_10198_), .C(_10647_), .Y(_10648_) );
	NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_10648_), .B(_10646_), .Y(_10649_) );
	AOI22X1 AOI22X1_572 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf2), .B(csr_gpr_iu_csr_sepc_22_), .C(csr_gpr_iu_csr_scause_22_), .D(_7435__bF_buf5), .Y(_10650_) );
	OAI21X1 OAI21X1_4324 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .B(_8617_), .C(_10650_), .Y(_10651_) );
	AOI22X1 AOI22X1_573 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_22_), .B(_8233__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_22_), .D(_8280__bF_buf4), .Y(_10652_) );
	AOI22X1 AOI22X1_574 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_22_), .B(_8846__bF_buf3), .C(csr_gpr_iu_csr_mscratch_22_), .D(_8417__bF_buf3), .Y(_10653_) );
	AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_10652_), .B(_10653_), .Y(_10654_) );
	OAI21X1 OAI21X1_4325 ( .gnd(gnd), .vdd(vdd), .A(_8795_), .B(_10215_), .C(_10654_), .Y(_10655_) );
	NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_10651_), .B(_10655_), .Y(_10656_) );
	NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(_10644_), .B(_10649_), .C(_10656_), .Y(csr_22_) );
	AOI22X1 AOI22X1_575 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_23_), .B(_8062__bF_buf1), .C(csr_gpr_iu_csr_mcycle_23_), .D(_10165_), .Y(_10657_) );
	OAI21X1 OAI21X1_4326 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_9161__bF_buf2), .C(_10657_), .Y(_10658_) );
	OAI21X1 OAI21X1_4327 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_23_), .B(csr_gpr_iu_csr_mideleg_23_), .C(_10170_), .Y(_10659_) );
	AOI22X1 AOI22X1_576 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_23_), .B(_10163_), .C(csr_gpr_iu_csr_minstret_23_), .D(_10227_), .Y(_10660_) );
	AOI22X1 AOI22X1_577 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf1), .B(csr_gpr_iu_csr_pmpaddr2_23_), .C(csr_gpr_iu_csr_mtval_23_), .D(_8618__bF_buf2), .Y(_10661_) );
	NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(_10659_), .B(_10661_), .C(_10660_), .Y(_10662_) );
	NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_10658_), .B(_10662_), .Y(_10663_) );
	OAI22X1 OAI22X1_802 ( .gnd(gnd), .vdd(vdd), .A(_8147_), .B(_8116_), .C(_8029_), .D(_7959_), .Y(_10664_) );
	OAI22X1 OAI22X1_803 ( .gnd(gnd), .vdd(vdd), .A(_8351_), .B(_8326_), .C(_8396_), .D(_8371_), .Y(_10665_) );
	NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_10665_), .B(_10664_), .Y(_10666_) );
	AOI22X1 AOI22X1_578 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf1), .B(csr_gpr_iu_csr_sepc_23_), .C(csr_gpr_iu_csr_mcause_23_), .D(_10235_), .Y(_10667_) );
	AOI22X1 AOI22X1_579 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf4), .B(csr_gpr_iu_csr_scause_23_), .C(csr_gpr_iu_csr_pmpaddr1_23_), .D(_8233__bF_buf2), .Y(_10668_) );
	NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_10668_), .B(_10667_), .Y(_10669_) );
	AOI22X1 AOI22X1_580 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_23_), .B(_8846__bF_buf2), .C(csr_gpr_iu_csr_mscratch_23_), .D(_8417__bF_buf2), .Y(_10670_) );
	AOI22X1 AOI22X1_581 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_23_), .B(_7323__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_23_), .D(_8280__bF_buf3), .Y(_10671_) );
	NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_10670_), .B(_10671_), .Y(_10672_) );
	NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_10669_), .B(_10672_), .Y(_10673_) );
	NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(_10666_), .B(_10673_), .C(_10663_), .Y(csr_23_) );
	OAI22X1 OAI22X1_804 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9019__bF_buf3), .C(_7236_), .D(_10164_), .Y(_10674_) );
	AOI21X1 AOI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_24_), .B(_10227_), .C(_10674_), .Y(_10675_) );
	AOI22X1 AOI22X1_582 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf2), .B(biu_mmu_satp_24_), .C(csr_gpr_iu_csr_stvec_24_), .D(_8062__bF_buf0), .Y(_10676_) );
	OAI21X1 OAI21X1_4328 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_8684__bF_buf5), .C(_10676_), .Y(_10677_) );
	OAI21X1 OAI21X1_4329 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_24_), .B(csr_gpr_iu_csr_mideleg_24_), .C(_10170_), .Y(_10678_) );
	OAI21X1 OAI21X1_4330 ( .gnd(gnd), .vdd(vdd), .A(_8032_), .B(_7959_), .C(_10678_), .Y(_10679_) );
	NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_10677_), .B(_10679_), .Y(_10680_) );
	AOI22X1 AOI22X1_583 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf0), .B(csr_gpr_iu_csr_sscratch_24_), .C(csr_gpr_iu_csr_sepc_24_), .D(_7584__bF_buf0), .Y(_10681_) );
	AOI22X1 AOI22X1_584 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_24_), .B(_8233__bF_buf1), .C(csr_gpr_iu_csr_mscratch_24_), .D(_8417__bF_buf1), .Y(_10682_) );
	NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_10681_), .B(_10682_), .Y(_10683_) );
	AOI22X1 AOI22X1_585 ( .gnd(gnd), .vdd(vdd), .A(_8280__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr0_24_), .C(csr_gpr_iu_csr_mtval_24_), .D(_8618__bF_buf1), .Y(_10684_) );
	AOI22X1 AOI22X1_586 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_24_), .B(_8846__bF_buf1), .C(csr_gpr_iu_csr_pmp3cfg_0_), .D(_8372__bF_buf5), .Y(_10685_) );
	AOI22X1 AOI22X1_587 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_24_), .B(_7435__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr3_24_), .D(_8117__bF_buf6), .Y(_10686_) );
	AOI22X1 AOI22X1_588 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_0_), .B(_8327__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr2_24_), .D(_10182__bF_buf0), .Y(_10687_) );
	AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_10686_), .B(_10687_), .Y(_10688_) );
	NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_10684_), .B(_10685_), .C(_10688_), .Y(_10689_) );
	NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_10683_), .B(_10689_), .Y(_10690_) );
	NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_10675_), .B(_10680_), .C(_10690_), .Y(csr_24_) );
	AOI22X1 AOI22X1_589 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_25_), .B(_8062__bF_buf5), .C(csr_gpr_iu_csr_mcycle_25_), .D(_10165_), .Y(_10691_) );
	OAI21X1 OAI21X1_4331 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_9161__bF_buf1), .C(_10691_), .Y(_10692_) );
	OAI21X1 OAI21X1_4332 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_25_), .B(csr_gpr_iu_csr_mideleg_25_), .C(_10170_), .Y(_10693_) );
	AOI22X1 AOI22X1_590 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_25_), .B(_10163_), .C(csr_gpr_iu_csr_minstret_25_), .D(_10227_), .Y(_10694_) );
	AOI22X1 AOI22X1_591 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf3), .B(csr_gpr_iu_csr_pmpaddr2_25_), .C(csr_gpr_iu_csr_mtval_25_), .D(_8618__bF_buf0), .Y(_10695_) );
	NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_10693_), .B(_10695_), .C(_10694_), .Y(_10696_) );
	NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_10692_), .B(_10696_), .Y(_10697_) );
	OAI22X1 OAI22X1_805 ( .gnd(gnd), .vdd(vdd), .A(_8150_), .B(_8116_), .C(_7543_), .D(_7437_), .Y(_10698_) );
	OAI22X1 OAI22X1_806 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(_8232_), .C(_8330_), .D(_8326_), .Y(_10699_) );
	NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_10699_), .B(_10698_), .Y(_10700_) );
	AOI22X1 AOI22X1_592 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf5), .B(csr_gpr_iu_csr_sepc_25_), .C(csr_gpr_iu_csr_mcause_25_), .D(_10235_), .Y(_10701_) );
	AOI22X1 AOI22X1_593 ( .gnd(gnd), .vdd(vdd), .A(_8280__bF_buf1), .B(csr_gpr_iu_csr_pmpaddr0_25_), .C(csr_gpr_iu_csr_pmp3cfg_1_), .D(_8372__bF_buf4), .Y(_10702_) );
	NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_10701_), .B(_10702_), .Y(_10703_) );
	AOI22X1 AOI22X1_594 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_25_), .B(_8846__bF_buf0), .C(csr_gpr_iu_csr_mscratch_25_), .D(_8417__bF_buf0), .Y(_10704_) );
	AOI22X1 AOI22X1_595 ( .gnd(gnd), .vdd(vdd), .A(_7323__bF_buf1), .B(csr_gpr_iu_csr_sscratch_25_), .C(csr_gpr_iu_csr_stval_25_), .D(_7960__bF_buf5), .Y(_10705_) );
	NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_10704_), .B(_10705_), .Y(_10706_) );
	NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_10703_), .B(_10706_), .Y(_10707_) );
	NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(_10700_), .B(_10697_), .C(_10707_), .Y(csr_25_) );
	AOI22X1 AOI22X1_596 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_26_), .B(_10163_), .C(csr_gpr_iu_csr_mcycle_26_), .D(_10165_), .Y(_10708_) );
	OAI21X1 OAI21X1_4333 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_10162_), .C(_10708_), .Y(_10709_) );
	NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_26_), .B(_9234__bF_buf1), .Y(_10710_) );
	OAI21X1 OAI21X1_4334 ( .gnd(gnd), .vdd(vdd), .A(_9999_), .B(_8061_), .C(_10710_), .Y(_10711_) );
	AOI21X1 AOI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcause_26_), .B(_10235_), .C(_10711_), .Y(_10712_) );
	NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stval_26_), .B(_7960__bF_buf4), .Y(_10713_) );
	OAI21X1 OAI21X1_4335 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_26_), .B(csr_gpr_iu_csr_mideleg_26_), .C(_10170_), .Y(_10714_) );
	NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10714_), .C(_10712_), .Y(_10715_) );
	NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .B(_10715_), .Y(_10716_) );
	AOI22X1 AOI22X1_597 ( .gnd(gnd), .vdd(vdd), .A(_7319__bF_buf4), .B(csr_gpr_iu_csr_sscratch_26_), .C(csr_gpr_iu_csr_sepc_26_), .D(_7584__bF_buf4), .Y(_10717_) );
	AOI22X1 AOI22X1_598 ( .gnd(gnd), .vdd(vdd), .A(_8280__bF_buf0), .B(csr_gpr_iu_csr_pmpaddr0_26_), .C(csr_gpr_iu_csr_mscratch_26_), .D(_8417__bF_buf5), .Y(_10718_) );
	AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_10718_), .B(_10717_), .Y(_10719_) );
	AOI22X1 AOI22X1_599 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_26_), .B(_8233__bF_buf0), .C(csr_gpr_iu_csr_mtval_26_), .D(_8618__bF_buf6), .Y(_10720_) );
	AOI22X1 AOI22X1_600 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_26_), .B(_8846__bF_buf3), .C(csr_gpr_iu_csr_pmp3cfg_2_), .D(_8372__bF_buf3), .Y(_10721_) );
	NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_10721_), .B(_10720_), .Y(_10722_) );
	NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_26_), .B(_8117__bF_buf5), .Y(_10723_) );
	NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_26_), .B(_7435__bF_buf2), .Y(_10724_) );
	AOI22X1 AOI22X1_601 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_2_), .B(_8327__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr2_26_), .D(_10182__bF_buf2), .Y(_10725_) );
	NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_10723_), .B(_10724_), .C(_10725_), .Y(_10726_) );
	NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_10722_), .B(_10726_), .Y(_10727_) );
	NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_10719_), .B(_10727_), .C(_10716_), .Y(csr_26_) );
	AOI22X1 AOI22X1_602 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mcycle_27_), .B(_10186_), .C(csr_gpr_iu_csr_minstret_27_), .D(_10208_), .Y(_10728_) );
	OAI21X1 OAI21X1_4336 ( .gnd(gnd), .vdd(vdd), .A(_9077_), .B(_9019__bF_buf2), .C(_10728_), .Y(_10729_) );
	AOI21X1 AOI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mscratch_27_), .B(_8417__bF_buf4), .C(_10729_), .Y(_10730_) );
	OAI22X1 OAI22X1_807 ( .gnd(gnd), .vdd(vdd), .A(_8674_), .B(_8617_), .C(_8820_), .D(_10215_), .Y(_10731_) );
	AOI21X1 AOI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_27_), .B(_8846__bF_buf2), .C(_10731_), .Y(_10732_) );
	NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_8544_), .B(_8602_), .Y(_10733_) );
	AOI22X1 AOI22X1_603 ( .gnd(gnd), .vdd(vdd), .A(_8165__bF_buf0), .B(csr_gpr_iu_csr_pmpaddr2_27_), .C(_8489__bF_buf3), .D(_10733_), .Y(_10734_) );
	NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(_10734_), .B(_10732_), .C(_10730_), .Y(_10735_) );
	OAI22X1 OAI22X1_808 ( .gnd(gnd), .vdd(vdd), .A(_7408_), .B(_7320__bF_buf0), .C(_7895_), .D(_7586__bF_buf3), .Y(_10736_) );
	AOI21X1 AOI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_27_), .B(_8062__bF_buf4), .C(_10736_), .Y(_10737_) );
	AOI22X1 AOI22X1_604 ( .gnd(gnd), .vdd(vdd), .A(_8117__bF_buf4), .B(csr_gpr_iu_csr_pmpaddr3_27_), .C(csr_gpr_iu_csr_pmp3cfg_3_), .D(_8372__bF_buf2), .Y(_10738_) );
	AOI22X1 AOI22X1_605 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf1), .B(csr_gpr_iu_csr_scause_27_), .C(csr_gpr_iu_csr_stval_27_), .D(_10199_), .Y(_10739_) );
	OAI21X1 OAI21X1_4337 ( .gnd(gnd), .vdd(vdd), .A(_9221_), .B(_9161__bF_buf0), .C(_10739_), .Y(_10740_) );
	AOI22X1 AOI22X1_606 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_27_), .B(_8233__bF_buf5), .C(csr_gpr_iu_csr_pmpaddr0_27_), .D(_8280__bF_buf5), .Y(_10741_) );
	OAI21X1 OAI21X1_4338 ( .gnd(gnd), .vdd(vdd), .A(_8333_), .B(_8326_), .C(_10741_), .Y(_10742_) );
	NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_10740_), .B(_10742_), .Y(_10743_) );
	NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .B(_10738_), .C(_10743_), .Y(_10744_) );
	OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_10744_), .B(_10735_), .Y(csr_27_) );
	OAI22X1 OAI22X1_809 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9019__bF_buf1), .C(_7259_), .D(_10164_), .Y(_10745_) );
	AOI21X1 AOI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_minstret_28_), .B(_10227_), .C(_10745_), .Y(_10746_) );
	AOI22X1 AOI22X1_607 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf0), .B(biu_mmu_satp_28_), .C(csr_gpr_iu_csr_stvec_28_), .D(_8062__bF_buf3), .Y(_10747_) );
	OAI21X1 OAI21X1_4339 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_8684__bF_buf4), .C(_10747_), .Y(_10748_) );
	INVX1 INVX1_1700 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr0_28_), .Y(_10749_) );
	OAI21X1 OAI21X1_4340 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_28_), .B(csr_gpr_iu_csr_mideleg_28_), .C(_10170_), .Y(_10750_) );
	OAI21X1 OAI21X1_4341 ( .gnd(gnd), .vdd(vdd), .A(_10749_), .B(_8279_), .C(_10750_), .Y(_10751_) );
	NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_10748_), .B(_10751_), .Y(_10752_) );
	NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sepc_28_), .B(_7584__bF_buf3), .Y(_10753_) );
	NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_28_), .B(_7323__bF_buf0), .Y(_10754_) );
	AOI22X1 AOI22X1_608 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr1_28_), .B(_8233__bF_buf4), .C(csr_gpr_iu_csr_mscratch_28_), .D(_8417__bF_buf3), .Y(_10755_) );
	NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .B(_10754_), .C(_10755_), .Y(_10756_) );
	NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_4_), .B(_8327__bF_buf1), .Y(_10757_) );
	OAI21X1 OAI21X1_4342 ( .gnd(gnd), .vdd(vdd), .A(_8676_), .B(_8617_), .C(_10757_), .Y(_10758_) );
	OAI22X1 OAI22X1_810 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8847__bF_buf2), .C(_7558_), .D(_7437_), .Y(_10759_) );
	NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_10759_), .B(_10758_), .Y(_10760_) );
	AOI22X1 AOI22X1_609 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_28_), .B(_8117__bF_buf3), .C(csr_gpr_iu_csr_stval_28_), .D(_7960__bF_buf3), .Y(_10761_) );
	AOI22X1 AOI22X1_610 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf1), .B(csr_gpr_iu_csr_pmpaddr2_28_), .C(csr_gpr_iu_csr_pmp3cfg_4_), .D(_8372__bF_buf1), .Y(_10762_) );
	NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_10761_), .B(_10762_), .C(_10760_), .Y(_10763_) );
	NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_10756_), .B(_10763_), .Y(_10764_) );
	NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(_10746_), .B(_10752_), .C(_10764_), .Y(csr_28_) );
	AOI22X1 AOI22X1_611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_29_), .B(_8062__bF_buf2), .C(csr_gpr_iu_csr_mcycle_29_), .D(_10165_), .Y(_10765_) );
	OAI21X1 OAI21X1_4343 ( .gnd(gnd), .vdd(vdd), .A(_9225_), .B(_9161__bF_buf4), .C(_10765_), .Y(_10766_) );
	OAI21X1 OAI21X1_4344 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_29_), .B(csr_gpr_iu_csr_mideleg_29_), .C(_10170_), .Y(_10767_) );
	AOI22X1 AOI22X1_612 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_29_), .B(_10163_), .C(csr_gpr_iu_csr_minstret_29_), .D(_10227_), .Y(_10768_) );
	AOI22X1 AOI22X1_613 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf0), .B(csr_gpr_iu_csr_pmpaddr2_29_), .C(csr_gpr_iu_csr_mtval_29_), .D(_8618__bF_buf5), .Y(_10769_) );
	NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(_10767_), .B(_10769_), .C(_10768_), .Y(_10770_) );
	NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10770_), .Y(_10771_) );
	AOI22X1 AOI22X1_614 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_29_), .B(_8117__bF_buf2), .C(csr_gpr_iu_csr_stval_29_), .D(_7960__bF_buf2), .Y(_10772_) );
	AOI22X1 AOI22X1_615 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_5_), .B(_8327__bF_buf0), .C(csr_gpr_iu_csr_pmp3cfg_5_), .D(_8372__bF_buf0), .Y(_10773_) );
	NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_10773_), .B(_10772_), .Y(_10774_) );
	OAI22X1 OAI22X1_811 ( .gnd(gnd), .vdd(vdd), .A(_8830_), .B(_8684__bF_buf3), .C(_7913_), .D(_7586__bF_buf2), .Y(_10775_) );
	NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_scause_29_), .B(_7435__bF_buf0), .Y(_10776_) );
	OAI21X1 OAI21X1_4345 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .B(_8232_), .C(_10776_), .Y(_10777_) );
	NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_10777_), .B(_10775_), .Y(_10778_) );
	AOI22X1 AOI22X1_616 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_29_), .B(_8846__bF_buf1), .C(csr_gpr_iu_csr_mscratch_29_), .D(_8417__bF_buf2), .Y(_10779_) );
	AOI22X1 AOI22X1_617 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_29_), .B(_7323__bF_buf3), .C(csr_gpr_iu_csr_pmpaddr0_29_), .D(_8280__bF_buf4), .Y(_10780_) );
	NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_10779_), .B(_10780_), .C(_10778_), .Y(_10781_) );
	NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_10774_), .B(_10781_), .Y(_10782_) );
	NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_10771_), .B(_10782_), .Y(csr_29_) );
	INVX1 INVX1_1701 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_satp_30_), .Y(_10783_) );
	AOI22X1 AOI22X1_618 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stvec_30_), .B(_8062__bF_buf1), .C(csr_gpr_iu_csr_mcycle_30_), .D(_10165_), .Y(_10784_) );
	OAI21X1 OAI21X1_4346 ( .gnd(gnd), .vdd(vdd), .A(_10783_), .B(_9161__bF_buf3), .C(_10784_), .Y(_10785_) );
	OAI21X1 OAI21X1_4347 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_30_), .B(csr_gpr_iu_csr_mideleg_30_), .C(_10170_), .Y(_10786_) );
	AOI22X1 AOI22X1_619 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_30_), .B(_10163_), .C(csr_gpr_iu_csr_minstret_30_), .D(_10227_), .Y(_10787_) );
	AOI22X1 AOI22X1_620 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf3), .B(csr_gpr_iu_csr_pmpaddr2_30_), .C(csr_gpr_iu_csr_mtval_30_), .D(_8618__bF_buf4), .Y(_10788_) );
	NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10788_), .C(_10787_), .Y(_10789_) );
	NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_10785_), .B(_10789_), .Y(_10790_) );
	AOI22X1 AOI22X1_621 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_30_), .B(_8117__bF_buf1), .C(csr_gpr_iu_csr_stval_30_), .D(_7960__bF_buf1), .Y(_10791_) );
	AOI22X1 AOI22X1_622 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_6_), .B(_8327__bF_buf6), .C(csr_gpr_iu_csr_pmp3cfg_6_), .D(_8372__bF_buf6), .Y(_10792_) );
	AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_10791_), .B(_10792_), .Y(_10793_) );
	AOI22X1 AOI22X1_623 ( .gnd(gnd), .vdd(vdd), .A(_7584__bF_buf2), .B(csr_gpr_iu_csr_sepc_30_), .C(csr_gpr_iu_csr_mcause_30_), .D(_10235_), .Y(_10794_) );
	AOI22X1 AOI22X1_624 ( .gnd(gnd), .vdd(vdd), .A(_7435__bF_buf6), .B(csr_gpr_iu_csr_scause_30_), .C(csr_gpr_iu_csr_pmpaddr1_30_), .D(_8233__bF_buf3), .Y(_10795_) );
	NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_10795_), .B(_10794_), .Y(_10796_) );
	AOI22X1 AOI22X1_625 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_30_), .B(_8846__bF_buf0), .C(csr_gpr_iu_csr_mscratch_30_), .D(_8417__bF_buf1), .Y(_10797_) );
	AOI22X1 AOI22X1_626 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sscratch_30_), .B(_7323__bF_buf2), .C(csr_gpr_iu_csr_pmpaddr0_30_), .D(_8280__bF_buf3), .Y(_10798_) );
	NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_10797_), .B(_10798_), .Y(_10799_) );
	NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .B(_10799_), .Y(_10800_) );
	NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_10793_), .B(_10800_), .C(_10790_), .Y(csr_30_) );
	AOI22X1 AOI22X1_627 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mtvec_31_), .B(_10163_), .C(csr_gpr_iu_csr_mcycle_31_), .D(_10165_), .Y(_10801_) );
	OAI21X1 OAI21X1_4348 ( .gnd(gnd), .vdd(vdd), .A(_6854_), .B(_10162_), .C(_10801_), .Y(_10802_) );
	AOI22X1 AOI22X1_628 ( .gnd(gnd), .vdd(vdd), .A(_9234__bF_buf3), .B(biu_mmu_satp_31_), .C(csr_gpr_iu_csr_stvec_31_), .D(_8062__bF_buf0), .Y(_10803_) );
	OAI21X1 OAI21X1_4349 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(_8684__bF_buf2), .C(_10803_), .Y(_10804_) );
	OAI21X1 OAI21X1_4350 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_31_), .B(csr_gpr_iu_csr_mideleg_31_), .C(_10170_), .Y(_10805_) );
	OAI21X1 OAI21X1_4351 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(_8279_), .C(_10805_), .Y(_10806_) );
	OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_10806_), .B(_10804_), .Y(_10807_) );
	NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_10802_), .B(_10807_), .Y(_10808_) );
	OAI22X1 OAI22X1_812 ( .gnd(gnd), .vdd(vdd), .A(_7948_), .B(_7586__bF_buf1), .C(_7419_), .D(_9233_), .Y(_10809_) );
	OAI22X1 OAI22X1_813 ( .gnd(gnd), .vdd(vdd), .A(_8276_), .B(_8232_), .C(_8464_), .D(_8416_), .Y(_10810_) );
	NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_10810_), .B(_10809_), .Y(_10811_) );
	AOI22X1 AOI22X1_629 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmp7cfg_7_), .B(_8327__bF_buf5), .C(csr_gpr_iu_csr_mtval_31_), .D(_8618__bF_buf3), .Y(_10812_) );
	AOI22X1 AOI22X1_630 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mepc_31_), .B(_8846__bF_buf3), .C(csr_gpr_iu_csr_scause_31_bF_buf1), .D(_7435__bF_buf5), .Y(_10813_) );
	NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_10813_), .B(_10812_), .Y(_10814_) );
	AOI22X1 AOI22X1_631 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pmpaddr3_31_), .B(_8117__bF_buf0), .C(csr_gpr_iu_csr_stval_31_), .D(_7960__bF_buf0), .Y(_10815_) );
	AOI22X1 AOI22X1_632 ( .gnd(gnd), .vdd(vdd), .A(_10182__bF_buf2), .B(csr_gpr_iu_csr_pmpaddr2_31_), .C(csr_gpr_iu_csr_pmp3cfg_7_), .D(_8372__bF_buf5), .Y(_10816_) );
	NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_10816_), .B(_10815_), .Y(_10817_) );
	NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_10814_), .B(_10817_), .Y(_10818_) );
	NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(_10811_), .B(_10818_), .C(_10808_), .Y(csr_31_) );
	DFFPOSX1 DFFPOSX1_1178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6705__0_), .Q(csr_gpr_iu_csr_mcycle_0_) );
	DFFPOSX1 DFFPOSX1_1179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6705__1_), .Q(csr_gpr_iu_csr_mcycle_1_) );
	DFFPOSX1 DFFPOSX1_1180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6705__2_), .Q(csr_gpr_iu_csr_mcycle_2_) );
	DFFPOSX1 DFFPOSX1_1181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6705__3_), .Q(csr_gpr_iu_csr_mcycle_3_) );
	DFFPOSX1 DFFPOSX1_1182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6705__4_), .Q(csr_gpr_iu_csr_mcycle_4_) );
	DFFPOSX1 DFFPOSX1_1183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6705__5_), .Q(csr_gpr_iu_csr_mcycle_5_) );
	DFFPOSX1 DFFPOSX1_1184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6705__6_), .Q(csr_gpr_iu_csr_mcycle_6_) );
	DFFPOSX1 DFFPOSX1_1185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6705__7_), .Q(csr_gpr_iu_csr_mcycle_7_) );
	DFFPOSX1 DFFPOSX1_1186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6705__8_), .Q(csr_gpr_iu_csr_mcycle_8_) );
	DFFPOSX1 DFFPOSX1_1187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6705__9_), .Q(csr_gpr_iu_csr_mcycle_9_) );
	DFFPOSX1 DFFPOSX1_1188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6705__10_), .Q(csr_gpr_iu_csr_mcycle_10_) );
	DFFPOSX1 DFFPOSX1_1189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6705__11_), .Q(csr_gpr_iu_csr_mcycle_11_) );
	DFFPOSX1 DFFPOSX1_1190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6705__12_), .Q(csr_gpr_iu_csr_mcycle_12_) );
	DFFPOSX1 DFFPOSX1_1191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6705__13_), .Q(csr_gpr_iu_csr_mcycle_13_) );
	DFFPOSX1 DFFPOSX1_1192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6705__14_), .Q(csr_gpr_iu_csr_mcycle_14_) );
	DFFPOSX1 DFFPOSX1_1193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_6705__15_), .Q(csr_gpr_iu_csr_mcycle_15_) );
	DFFPOSX1 DFFPOSX1_1194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_6705__16_), .Q(csr_gpr_iu_csr_mcycle_16_) );
	DFFPOSX1 DFFPOSX1_1195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_6705__17_), .Q(csr_gpr_iu_csr_mcycle_17_) );
	DFFPOSX1 DFFPOSX1_1196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_6705__18_), .Q(csr_gpr_iu_csr_mcycle_18_) );
	DFFPOSX1 DFFPOSX1_1197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_6705__19_), .Q(csr_gpr_iu_csr_mcycle_19_) );
	DFFPOSX1 DFFPOSX1_1198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_6705__20_), .Q(csr_gpr_iu_csr_mcycle_20_) );
	DFFPOSX1 DFFPOSX1_1199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_6705__21_), .Q(csr_gpr_iu_csr_mcycle_21_) );
	DFFPOSX1 DFFPOSX1_1200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_6705__22_), .Q(csr_gpr_iu_csr_mcycle_22_) );
	DFFPOSX1 DFFPOSX1_1201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_6705__23_), .Q(csr_gpr_iu_csr_mcycle_23_) );
	DFFPOSX1 DFFPOSX1_1202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_6705__24_), .Q(csr_gpr_iu_csr_mcycle_24_) );
	DFFPOSX1 DFFPOSX1_1203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_6705__25_), .Q(csr_gpr_iu_csr_mcycle_25_) );
	DFFPOSX1 DFFPOSX1_1204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_6705__26_), .Q(csr_gpr_iu_csr_mcycle_26_) );
	DFFPOSX1 DFFPOSX1_1205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_6705__27_), .Q(csr_gpr_iu_csr_mcycle_27_) );
	DFFPOSX1 DFFPOSX1_1206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_6705__28_), .Q(csr_gpr_iu_csr_mcycle_28_) );
	DFFPOSX1 DFFPOSX1_1207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_6705__29_), .Q(csr_gpr_iu_csr_mcycle_29_) );
	DFFPOSX1 DFFPOSX1_1208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_6705__30_), .Q(csr_gpr_iu_csr_mcycle_30_) );
	DFFPOSX1 DFFPOSX1_1209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_6705__31_), .Q(csr_gpr_iu_csr_mcycle_31_) );
	DFFPOSX1 DFFPOSX1_1210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_6712__0_), .Q(csr_gpr_iu_csr_minstret_0_) );
	DFFPOSX1 DFFPOSX1_1211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_6712__1_), .Q(csr_gpr_iu_csr_minstret_1_) );
	DFFPOSX1 DFFPOSX1_1212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_6712__2_), .Q(csr_gpr_iu_csr_minstret_2_) );
	DFFPOSX1 DFFPOSX1_1213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_6712__3_), .Q(csr_gpr_iu_csr_minstret_3_) );
	DFFPOSX1 DFFPOSX1_1214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_6712__4_), .Q(csr_gpr_iu_csr_minstret_4_) );
	DFFPOSX1 DFFPOSX1_1215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_6712__5_), .Q(csr_gpr_iu_csr_minstret_5_) );
	DFFPOSX1 DFFPOSX1_1216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_6712__6_), .Q(csr_gpr_iu_csr_minstret_6_) );
	DFFPOSX1 DFFPOSX1_1217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_6712__7_), .Q(csr_gpr_iu_csr_minstret_7_) );
	DFFPOSX1 DFFPOSX1_1218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_6712__8_), .Q(csr_gpr_iu_csr_minstret_8_) );
	DFFPOSX1 DFFPOSX1_1219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_6712__9_), .Q(csr_gpr_iu_csr_minstret_9_) );
	DFFPOSX1 DFFPOSX1_1220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_6712__10_), .Q(csr_gpr_iu_csr_minstret_10_) );
	DFFPOSX1 DFFPOSX1_1221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6712__11_), .Q(csr_gpr_iu_csr_minstret_11_) );
	DFFPOSX1 DFFPOSX1_1222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6712__12_), .Q(csr_gpr_iu_csr_minstret_12_) );
	DFFPOSX1 DFFPOSX1_1223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6712__13_), .Q(csr_gpr_iu_csr_minstret_13_) );
	DFFPOSX1 DFFPOSX1_1224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6712__14_), .Q(csr_gpr_iu_csr_minstret_14_) );
	DFFPOSX1 DFFPOSX1_1225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6712__15_), .Q(csr_gpr_iu_csr_minstret_15_) );
	DFFPOSX1 DFFPOSX1_1226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6712__16_), .Q(csr_gpr_iu_csr_minstret_16_) );
	DFFPOSX1 DFFPOSX1_1227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6712__17_), .Q(csr_gpr_iu_csr_minstret_17_) );
	DFFPOSX1 DFFPOSX1_1228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6712__18_), .Q(csr_gpr_iu_csr_minstret_18_) );
	DFFPOSX1 DFFPOSX1_1229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6712__19_), .Q(csr_gpr_iu_csr_minstret_19_) );
	DFFPOSX1 DFFPOSX1_1230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6712__20_), .Q(csr_gpr_iu_csr_minstret_20_) );
	DFFPOSX1 DFFPOSX1_1231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6712__21_), .Q(csr_gpr_iu_csr_minstret_21_) );
	DFFPOSX1 DFFPOSX1_1232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6712__22_), .Q(csr_gpr_iu_csr_minstret_22_) );
	DFFPOSX1 DFFPOSX1_1233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6712__23_), .Q(csr_gpr_iu_csr_minstret_23_) );
	DFFPOSX1 DFFPOSX1_1234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6712__24_), .Q(csr_gpr_iu_csr_minstret_24_) );
	DFFPOSX1 DFFPOSX1_1235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6712__25_), .Q(csr_gpr_iu_csr_minstret_25_) );
	DFFPOSX1 DFFPOSX1_1236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6712__26_), .Q(csr_gpr_iu_csr_minstret_26_) );
	DFFPOSX1 DFFPOSX1_1237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6712__27_), .Q(csr_gpr_iu_csr_minstret_27_) );
	DFFPOSX1 DFFPOSX1_1238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6712__28_), .Q(csr_gpr_iu_csr_minstret_28_) );
	DFFPOSX1 DFFPOSX1_1239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6712__29_), .Q(csr_gpr_iu_csr_minstret_29_) );
	DFFPOSX1 DFFPOSX1_1240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6712__30_), .Q(csr_gpr_iu_csr_minstret_30_) );
	DFFPOSX1 DFFPOSX1_1241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6712__31_), .Q(csr_gpr_iu_csr_minstret_31_) );
	DFFPOSX1 DFFPOSX1_1242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6708_), .Q(csr_gpr_iu_csr_meip) );
	DFFPOSX1 DFFPOSX1_1243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6741_), .Q(csr_gpr_iu_csr_seip) );
	DFFPOSX1 DFFPOSX1_1244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6721_), .Q(csr_gpr_iu_csr_mtip) );
	DFFPOSX1 DFFPOSX1_1245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6750_), .Q(csr_gpr_iu_csr_stip) );
	DFFPOSX1 DFFPOSX1_1246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6718_), .Q(csr_gpr_iu_csr_msip) );
	DFFPOSX1 DFFPOSX1_1247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6748_), .Q(csr_gpr_iu_csr_ssip) );
	DFFPOSX1 DFFPOSX1_1248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6725__0_), .Q(biu_pc_0_) );
	DFFPOSX1 DFFPOSX1_1249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6725__1_), .Q(biu_pc_1_) );
	DFFPOSX1 DFFPOSX1_1250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6725__2_), .Q(biu_pc_2_) );
	DFFPOSX1 DFFPOSX1_1251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6725__3_), .Q(biu_pc_3_) );
	DFFPOSX1 DFFPOSX1_1252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6725__4_), .Q(biu_pc_4_) );
	DFFPOSX1 DFFPOSX1_1253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6725__5_), .Q(biu_pc_5_) );
	DFFPOSX1 DFFPOSX1_1254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_6725__6_), .Q(biu_pc_6_) );
	DFFPOSX1 DFFPOSX1_1255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_6725__7_), .Q(biu_pc_7_) );
	DFFPOSX1 DFFPOSX1_1256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_6725__8_), .Q(biu_pc_8_) );
	DFFPOSX1 DFFPOSX1_1257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_6725__9_), .Q(biu_pc_9_) );
	DFFPOSX1 DFFPOSX1_1258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_6725__10_), .Q(biu_pc_10_) );
	DFFPOSX1 DFFPOSX1_1259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_6725__11_), .Q(biu_pc_11_) );
	DFFPOSX1 DFFPOSX1_1260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_6725__12_), .Q(biu_pc_12_) );
	DFFPOSX1 DFFPOSX1_1261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_6725__13_), .Q(biu_pc_13_) );
	DFFPOSX1 DFFPOSX1_1262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_6725__14_), .Q(biu_pc_14_) );
	DFFPOSX1 DFFPOSX1_1263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_6725__15_), .Q(biu_pc_15_) );
	DFFPOSX1 DFFPOSX1_1264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_6725__16_), .Q(biu_pc_16_) );
	DFFPOSX1 DFFPOSX1_1265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_6725__17_), .Q(biu_pc_17_) );
	DFFPOSX1 DFFPOSX1_1266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_6725__18_), .Q(biu_pc_18_) );
	DFFPOSX1 DFFPOSX1_1267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_6725__19_), .Q(biu_pc_19_) );
	DFFPOSX1 DFFPOSX1_1268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_6725__20_), .Q(biu_pc_20_) );
	DFFPOSX1 DFFPOSX1_1269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_6725__21_), .Q(biu_pc_21_) );
	DFFPOSX1 DFFPOSX1_1270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6725__22_), .Q(biu_pc_22_) );
	DFFPOSX1 DFFPOSX1_1271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_6725__23_), .Q(biu_pc_23_) );
	DFFPOSX1 DFFPOSX1_1272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_6725__24_), .Q(biu_pc_24_) );
	DFFPOSX1 DFFPOSX1_1273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_6725__25_), .Q(biu_pc_25_) );
	DFFPOSX1 DFFPOSX1_1274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_6725__26_), .Q(biu_pc_26_) );
	DFFPOSX1 DFFPOSX1_1275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_6725__27_), .Q(biu_pc_27_) );
	DFFPOSX1 DFFPOSX1_1276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_6725__28_), .Q(biu_pc_28_) );
	DFFPOSX1 DFFPOSX1_1277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_6725__29_), .Q(biu_pc_29_) );
	DFFPOSX1 DFFPOSX1_1278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6725__30_), .Q(biu_pc_30_) );
	DFFPOSX1 DFFPOSX1_1279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_6725__31_), .Q(biu_pc_31_) );
	DFFPOSX1 DFFPOSX1_1280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_6738__0_), .Q(biu_mmu_ag0_12_) );
	DFFPOSX1 DFFPOSX1_1281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_6738__1_), .Q(biu_mmu_ag0_13_) );
	DFFPOSX1 DFFPOSX1_1282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_6738__2_), .Q(biu_mmu_ag0_14_) );
	DFFPOSX1 DFFPOSX1_1283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_6738__3_), .Q(biu_mmu_ag0_15_) );
	DFFPOSX1 DFFPOSX1_1284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6738__4_), .Q(biu_mmu_ag0_16_) );
	DFFPOSX1 DFFPOSX1_1285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6738__5_), .Q(biu_mmu_ag0_17_) );
	DFFPOSX1 DFFPOSX1_1286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_6738__6_), .Q(biu_mmu_ag0_18_) );
	DFFPOSX1 DFFPOSX1_1287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6738__7_), .Q(biu_mmu_ag0_19_) );
	DFFPOSX1 DFFPOSX1_1288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6738__8_), .Q(biu_mmu_ag0_20_) );
	DFFPOSX1 DFFPOSX1_1289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_6738__9_), .Q(biu_mmu_ag0_21_) );
	DFFPOSX1 DFFPOSX1_1290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_6738__10_), .Q(biu_mmu_ag0_22_) );
	DFFPOSX1 DFFPOSX1_1291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_6738__11_), .Q(biu_mmu_ag0_23_) );
	DFFPOSX1 DFFPOSX1_1292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_6738__12_), .Q(biu_mmu_ag0_24_) );
	DFFPOSX1 DFFPOSX1_1293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_6738__13_), .Q(biu_mmu_ag0_25_) );
	DFFPOSX1 DFFPOSX1_1294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_6738__14_), .Q(biu_mmu_ag0_26_) );
	DFFPOSX1 DFFPOSX1_1295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_6738__15_), .Q(biu_mmu_ag0_27_) );
	DFFPOSX1 DFFPOSX1_1296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_6738__16_), .Q(biu_mmu_ag0_28_) );
	DFFPOSX1 DFFPOSX1_1297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_6738__17_), .Q(biu_mmu_ag0_29_) );
	DFFPOSX1 DFFPOSX1_1298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_6738__18_), .Q(biu_mmu_ag0_30_) );
	DFFPOSX1 DFFPOSX1_1299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_6738__19_), .Q(biu_mmu_ag0_31_) );
	DFFPOSX1 DFFPOSX1_1300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_6738__20_), .Q(biu_mmu_ag0_32_) );
	DFFPOSX1 DFFPOSX1_1301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_6738__21_), .Q(biu_mmu_ag0_33_) );
	DFFPOSX1 DFFPOSX1_1302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_6738__22_), .Q(biu_mmu_satp_22_) );
	DFFPOSX1 DFFPOSX1_1303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_6738__23_), .Q(biu_mmu_satp_23_) );
	DFFPOSX1 DFFPOSX1_1304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_6738__24_), .Q(biu_mmu_satp_24_) );
	DFFPOSX1 DFFPOSX1_1305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_6738__25_), .Q(biu_mmu_satp_25_) );
	DFFPOSX1 DFFPOSX1_1306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_6738__26_), .Q(biu_mmu_satp_26_) );
	DFFPOSX1 DFFPOSX1_1307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_6738__27_), .Q(biu_mmu_satp_27_) );
	DFFPOSX1 DFFPOSX1_1308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_6738__28_), .Q(biu_mmu_satp_28_) );
	DFFPOSX1 DFFPOSX1_1309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_6738__29_), .Q(biu_mmu_satp_29_) );
	DFFPOSX1 DFFPOSX1_1310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_6738__30_), .Q(biu_mmu_satp_30_) );
	DFFPOSX1 DFFPOSX1_1311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_6738__31_), .Q(biu_mmu_satp_31_) );
	DFFPOSX1 DFFPOSX1_1312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_6719__0_), .Q(biu_mmu_msu_0_) );
	DFFPOSX1 DFFPOSX1_1313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_6719__1_), .Q(biu_mmu_msu_1_) );
	DFFPOSX1 DFFPOSX1_1314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_6724_), .Q(biu_mmu_mxr) );
	DFFPOSX1 DFFPOSX1_1315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_6753_), .Q(biu_mmu_sum) );
	DFFPOSX1 DFFPOSX1_1316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_6754_), .Q(csr_gpr_iu_csr_tsr) );
	DFFPOSX1 DFFPOSX1_1317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_6755_), .Q(csr_gpr_iu_csr_tvm) );
	DFFPOSX1 DFFPOSX1_1318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_6715_), .Q(csr_gpr_iu_csr_mprv) );
	DFFPOSX1 DFFPOSX1_1319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_6714__0_), .Q(csr_gpr_iu_csr_mpp_0_) );
	DFFPOSX1 DFFPOSX1_1320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_6714__1_), .Q(csr_gpr_iu_csr_mpp_1_) );
	DFFPOSX1 DFFPOSX1_1321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_6745_), .Q(csr_gpr_iu_csr_spp) );
	DFFPOSX1 DFFPOSX1_1322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_6713_), .Q(csr_gpr_iu_csr_mpie) );
	DFFPOSX1 DFFPOSX1_1323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_6744_), .Q(csr_gpr_iu_csr_spie) );
	DFFPOSX1 DFFPOSX1_1324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_6711_), .Q(csr_gpr_iu_csr_mie) );
	DFFPOSX1 DFFPOSX1_1325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_6743_), .Q(csr_gpr_iu_csr_sie) );
	DFFPOSX1 DFFPOSX1_1326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_6723__0_), .Q(csr_gpr_iu_csr_mtvec_0_) );
	DFFPOSX1 DFFPOSX1_1327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_6723__1_), .Q(csr_gpr_iu_csr_mtvec_1_) );
	DFFPOSX1 DFFPOSX1_1328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_6723__2_), .Q(csr_gpr_iu_csr_mtvec_2_) );
	DFFPOSX1 DFFPOSX1_1329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_6723__3_), .Q(csr_gpr_iu_csr_mtvec_3_) );
	DFFPOSX1 DFFPOSX1_1330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_6723__4_), .Q(csr_gpr_iu_csr_mtvec_4_) );
	DFFPOSX1 DFFPOSX1_1331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_6723__5_), .Q(csr_gpr_iu_csr_mtvec_5_) );
	DFFPOSX1 DFFPOSX1_1332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_6723__6_), .Q(csr_gpr_iu_csr_mtvec_6_) );
	DFFPOSX1 DFFPOSX1_1333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_6723__7_), .Q(csr_gpr_iu_csr_mtvec_7_) );
	DFFPOSX1 DFFPOSX1_1334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_6723__8_), .Q(csr_gpr_iu_csr_mtvec_8_) );
	DFFPOSX1 DFFPOSX1_1335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_6723__9_), .Q(csr_gpr_iu_csr_mtvec_9_) );
	DFFPOSX1 DFFPOSX1_1336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_6723__10_), .Q(csr_gpr_iu_csr_mtvec_10_) );
	DFFPOSX1 DFFPOSX1_1337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_6723__11_), .Q(csr_gpr_iu_csr_mtvec_11_) );
	DFFPOSX1 DFFPOSX1_1338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_6723__12_), .Q(csr_gpr_iu_csr_mtvec_12_) );
	DFFPOSX1 DFFPOSX1_1339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6723__13_), .Q(csr_gpr_iu_csr_mtvec_13_) );
	DFFPOSX1 DFFPOSX1_1340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6723__14_), .Q(csr_gpr_iu_csr_mtvec_14_) );
	DFFPOSX1 DFFPOSX1_1341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6723__15_), .Q(csr_gpr_iu_csr_mtvec_15_) );
	DFFPOSX1 DFFPOSX1_1342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6723__16_), .Q(csr_gpr_iu_csr_mtvec_16_) );
	DFFPOSX1 DFFPOSX1_1343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6723__17_), .Q(csr_gpr_iu_csr_mtvec_17_) );
	DFFPOSX1 DFFPOSX1_1344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6723__18_), .Q(csr_gpr_iu_csr_mtvec_18_) );
	DFFPOSX1 DFFPOSX1_1345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6723__19_), .Q(csr_gpr_iu_csr_mtvec_19_) );
	DFFPOSX1 DFFPOSX1_1346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6723__20_), .Q(csr_gpr_iu_csr_mtvec_20_) );
	DFFPOSX1 DFFPOSX1_1347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6723__21_), .Q(csr_gpr_iu_csr_mtvec_21_) );
	DFFPOSX1 DFFPOSX1_1348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6723__22_), .Q(csr_gpr_iu_csr_mtvec_22_) );
	DFFPOSX1 DFFPOSX1_1349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6723__23_), .Q(csr_gpr_iu_csr_mtvec_23_) );
	DFFPOSX1 DFFPOSX1_1350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6723__24_), .Q(csr_gpr_iu_csr_mtvec_24_) );
	DFFPOSX1 DFFPOSX1_1351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6723__25_), .Q(csr_gpr_iu_csr_mtvec_25_) );
	DFFPOSX1 DFFPOSX1_1352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6723__26_), .Q(csr_gpr_iu_csr_mtvec_26_) );
	DFFPOSX1 DFFPOSX1_1353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6723__27_), .Q(csr_gpr_iu_csr_mtvec_27_) );
	DFFPOSX1 DFFPOSX1_1354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_6723__28_), .Q(csr_gpr_iu_csr_mtvec_28_) );
	DFFPOSX1 DFFPOSX1_1355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_6723__29_), .Q(csr_gpr_iu_csr_mtvec_29_) );
	DFFPOSX1 DFFPOSX1_1356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_6723__30_), .Q(csr_gpr_iu_csr_mtvec_30_) );
	DFFPOSX1 DFFPOSX1_1357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_6723__31_), .Q(csr_gpr_iu_csr_mtvec_31_) );
	DFFPOSX1 DFFPOSX1_1358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_6709__0_), .Q(csr_gpr_iu_csr_mepc_0_) );
	DFFPOSX1 DFFPOSX1_1359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_6709__1_), .Q(csr_gpr_iu_csr_mepc_1_) );
	DFFPOSX1 DFFPOSX1_1360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_6709__2_), .Q(csr_gpr_iu_csr_mepc_2_) );
	DFFPOSX1 DFFPOSX1_1361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_6709__3_), .Q(csr_gpr_iu_csr_mepc_3_) );
	DFFPOSX1 DFFPOSX1_1362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_6709__4_), .Q(csr_gpr_iu_csr_mepc_4_) );
	DFFPOSX1 DFFPOSX1_1363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_6709__5_), .Q(csr_gpr_iu_csr_mepc_5_) );
	DFFPOSX1 DFFPOSX1_1364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_6709__6_), .Q(csr_gpr_iu_csr_mepc_6_) );
	DFFPOSX1 DFFPOSX1_1365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_6709__7_), .Q(csr_gpr_iu_csr_mepc_7_) );
	DFFPOSX1 DFFPOSX1_1366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_6709__8_), .Q(csr_gpr_iu_csr_mepc_8_) );
	DFFPOSX1 DFFPOSX1_1367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_6709__9_), .Q(csr_gpr_iu_csr_mepc_9_) );
	DFFPOSX1 DFFPOSX1_1368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_6709__10_), .Q(csr_gpr_iu_csr_mepc_10_) );
	DFFPOSX1 DFFPOSX1_1369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_6709__11_), .Q(csr_gpr_iu_csr_mepc_11_) );
	DFFPOSX1 DFFPOSX1_1370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_6709__12_), .Q(csr_gpr_iu_csr_mepc_12_) );
	DFFPOSX1 DFFPOSX1_1371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_6709__13_), .Q(csr_gpr_iu_csr_mepc_13_) );
	DFFPOSX1 DFFPOSX1_1372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_6709__14_), .Q(csr_gpr_iu_csr_mepc_14_) );
	DFFPOSX1 DFFPOSX1_1373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_6709__15_), .Q(csr_gpr_iu_csr_mepc_15_) );
	DFFPOSX1 DFFPOSX1_1374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_6709__16_), .Q(csr_gpr_iu_csr_mepc_16_) );
	DFFPOSX1 DFFPOSX1_1375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_6709__17_), .Q(csr_gpr_iu_csr_mepc_17_) );
	DFFPOSX1 DFFPOSX1_1376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_6709__18_), .Q(csr_gpr_iu_csr_mepc_18_) );
	DFFPOSX1 DFFPOSX1_1377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_6709__19_), .Q(csr_gpr_iu_csr_mepc_19_) );
	DFFPOSX1 DFFPOSX1_1378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_6709__20_), .Q(csr_gpr_iu_csr_mepc_20_) );
	DFFPOSX1 DFFPOSX1_1379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_6709__21_), .Q(csr_gpr_iu_csr_mepc_21_) );
	DFFPOSX1 DFFPOSX1_1380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_6709__22_), .Q(csr_gpr_iu_csr_mepc_22_) );
	DFFPOSX1 DFFPOSX1_1381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_6709__23_), .Q(csr_gpr_iu_csr_mepc_23_) );
	DFFPOSX1 DFFPOSX1_1382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6709__24_), .Q(csr_gpr_iu_csr_mepc_24_) );
	DFFPOSX1 DFFPOSX1_1383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6709__25_), .Q(csr_gpr_iu_csr_mepc_25_) );
	DFFPOSX1 DFFPOSX1_1384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6709__26_), .Q(csr_gpr_iu_csr_mepc_26_) );
	DFFPOSX1 DFFPOSX1_1385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6709__27_), .Q(csr_gpr_iu_csr_mepc_27_) );
	DFFPOSX1 DFFPOSX1_1386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6709__28_), .Q(csr_gpr_iu_csr_mepc_28_) );
	DFFPOSX1 DFFPOSX1_1387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6709__29_), .Q(csr_gpr_iu_csr_mepc_29_) );
	DFFPOSX1 DFFPOSX1_1388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6709__30_), .Q(csr_gpr_iu_csr_mepc_30_) );
	DFFPOSX1 DFFPOSX1_1389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6709__31_), .Q(csr_gpr_iu_csr_mepc_31_) );
	DFFPOSX1 DFFPOSX1_1390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6704__0_), .Q(csr_gpr_iu_csr_mcause_0_) );
	DFFPOSX1 DFFPOSX1_1391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6704__1_), .Q(csr_gpr_iu_csr_mcause_1_) );
	DFFPOSX1 DFFPOSX1_1392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6704__2_), .Q(csr_gpr_iu_csr_mcause_2_) );
	DFFPOSX1 DFFPOSX1_1393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6704__3_), .Q(csr_gpr_iu_csr_mcause_3_) );
	DFFPOSX1 DFFPOSX1_1394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6704__4_), .Q(csr_gpr_iu_csr_mcause_4_) );
	DFFPOSX1 DFFPOSX1_1395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6704__5_), .Q(csr_gpr_iu_csr_mcause_5_) );
	DFFPOSX1 DFFPOSX1_1396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6704__6_), .Q(csr_gpr_iu_csr_mcause_6_) );
	DFFPOSX1 DFFPOSX1_1397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6704__7_), .Q(csr_gpr_iu_csr_mcause_7_) );
	DFFPOSX1 DFFPOSX1_1398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6704__8_), .Q(csr_gpr_iu_csr_mcause_8_) );
	DFFPOSX1 DFFPOSX1_1399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6704__9_), .Q(csr_gpr_iu_csr_mcause_9_) );
	DFFPOSX1 DFFPOSX1_1400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6704__10_), .Q(csr_gpr_iu_csr_mcause_10_) );
	DFFPOSX1 DFFPOSX1_1401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6704__11_), .Q(csr_gpr_iu_csr_mcause_11_) );
	DFFPOSX1 DFFPOSX1_1402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6704__12_), .Q(csr_gpr_iu_csr_mcause_12_) );
	DFFPOSX1 DFFPOSX1_1403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6704__13_), .Q(csr_gpr_iu_csr_mcause_13_) );
	DFFPOSX1 DFFPOSX1_1404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6704__14_), .Q(csr_gpr_iu_csr_mcause_14_) );
	DFFPOSX1 DFFPOSX1_1405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6704__15_), .Q(csr_gpr_iu_csr_mcause_15_) );
	DFFPOSX1 DFFPOSX1_1406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6704__16_), .Q(csr_gpr_iu_csr_mcause_16_) );
	DFFPOSX1 DFFPOSX1_1407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6704__17_), .Q(csr_gpr_iu_csr_mcause_17_) );
	DFFPOSX1 DFFPOSX1_1408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6704__18_), .Q(csr_gpr_iu_csr_mcause_18_) );
	DFFPOSX1 DFFPOSX1_1409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6704__19_), .Q(csr_gpr_iu_csr_mcause_19_) );
	DFFPOSX1 DFFPOSX1_1410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6704__20_), .Q(csr_gpr_iu_csr_mcause_20_) );
	DFFPOSX1 DFFPOSX1_1411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6704__21_), .Q(csr_gpr_iu_csr_mcause_21_) );
	DFFPOSX1 DFFPOSX1_1412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6704__22_), .Q(csr_gpr_iu_csr_mcause_22_) );
	DFFPOSX1 DFFPOSX1_1413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6704__23_), .Q(csr_gpr_iu_csr_mcause_23_) );
	DFFPOSX1 DFFPOSX1_1414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6704__24_), .Q(csr_gpr_iu_csr_mcause_24_) );
	DFFPOSX1 DFFPOSX1_1415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_6704__25_), .Q(csr_gpr_iu_csr_mcause_25_) );
	DFFPOSX1 DFFPOSX1_1416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_6704__26_), .Q(csr_gpr_iu_csr_mcause_26_) );
	DFFPOSX1 DFFPOSX1_1417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_6704__27_), .Q(csr_gpr_iu_csr_mcause_27_) );
	DFFPOSX1 DFFPOSX1_1418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_6704__28_), .Q(csr_gpr_iu_csr_mcause_28_) );
	DFFPOSX1 DFFPOSX1_1419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_6704__29_), .Q(csr_gpr_iu_csr_mcause_29_) );
	DFFPOSX1 DFFPOSX1_1420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_6704__30_), .Q(csr_gpr_iu_csr_mcause_30_) );
	DFFPOSX1 DFFPOSX1_1421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_6704__31_), .Q(csr_gpr_iu_csr_mcause_31_) );
	DFFPOSX1 DFFPOSX1_1422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_6722__0_), .Q(csr_gpr_iu_csr_mtval_0_) );
	DFFPOSX1 DFFPOSX1_1423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_6722__1_), .Q(csr_gpr_iu_csr_mtval_1_) );
	DFFPOSX1 DFFPOSX1_1424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_6722__2_), .Q(csr_gpr_iu_csr_mtval_2_) );
	DFFPOSX1 DFFPOSX1_1425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_6722__3_), .Q(csr_gpr_iu_csr_mtval_3_) );
	DFFPOSX1 DFFPOSX1_1426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_6722__4_), .Q(csr_gpr_iu_csr_mtval_4_) );
	DFFPOSX1 DFFPOSX1_1427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_6722__5_), .Q(csr_gpr_iu_csr_mtval_5_) );
	DFFPOSX1 DFFPOSX1_1428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_6722__6_), .Q(csr_gpr_iu_csr_mtval_6_) );
	DFFPOSX1 DFFPOSX1_1429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_6722__7_), .Q(csr_gpr_iu_csr_mtval_7_) );
	DFFPOSX1 DFFPOSX1_1430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_6722__8_), .Q(csr_gpr_iu_csr_mtval_8_) );
	DFFPOSX1 DFFPOSX1_1431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6722__9_), .Q(csr_gpr_iu_csr_mtval_9_) );
	DFFPOSX1 DFFPOSX1_1432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_6722__10_), .Q(csr_gpr_iu_csr_mtval_10_) );
	DFFPOSX1 DFFPOSX1_1433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_6722__11_), .Q(csr_gpr_iu_csr_mtval_11_) );
	DFFPOSX1 DFFPOSX1_1434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_6722__12_), .Q(csr_gpr_iu_csr_mtval_12_) );
	DFFPOSX1 DFFPOSX1_1435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_6722__13_), .Q(csr_gpr_iu_csr_mtval_13_) );
	DFFPOSX1 DFFPOSX1_1436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_6722__14_), .Q(csr_gpr_iu_csr_mtval_14_) );
	DFFPOSX1 DFFPOSX1_1437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_6722__15_), .Q(csr_gpr_iu_csr_mtval_15_) );
	DFFPOSX1 DFFPOSX1_1438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_6722__16_), .Q(csr_gpr_iu_csr_mtval_16_) );
	DFFPOSX1 DFFPOSX1_1439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6722__17_), .Q(csr_gpr_iu_csr_mtval_17_) );
	DFFPOSX1 DFFPOSX1_1440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_6722__18_), .Q(csr_gpr_iu_csr_mtval_18_) );
	DFFPOSX1 DFFPOSX1_1441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_6722__19_), .Q(csr_gpr_iu_csr_mtval_19_) );
	DFFPOSX1 DFFPOSX1_1442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_6722__20_), .Q(csr_gpr_iu_csr_mtval_20_) );
	DFFPOSX1 DFFPOSX1_1443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_6722__21_), .Q(csr_gpr_iu_csr_mtval_21_) );
	DFFPOSX1 DFFPOSX1_1444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_6722__22_), .Q(csr_gpr_iu_csr_mtval_22_) );
	DFFPOSX1 DFFPOSX1_1445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6722__23_), .Q(csr_gpr_iu_csr_mtval_23_) );
	DFFPOSX1 DFFPOSX1_1446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6722__24_), .Q(csr_gpr_iu_csr_mtval_24_) );
	DFFPOSX1 DFFPOSX1_1447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_6722__25_), .Q(csr_gpr_iu_csr_mtval_25_) );
	DFFPOSX1 DFFPOSX1_1448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6722__26_), .Q(csr_gpr_iu_csr_mtval_26_) );
	DFFPOSX1 DFFPOSX1_1449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6722__27_), .Q(csr_gpr_iu_csr_mtval_27_) );
	DFFPOSX1 DFFPOSX1_1450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_6722__28_), .Q(csr_gpr_iu_csr_mtval_28_) );
	DFFPOSX1 DFFPOSX1_1451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_6722__29_), .Q(csr_gpr_iu_csr_mtval_29_) );
	DFFPOSX1 DFFPOSX1_1452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_6722__30_), .Q(csr_gpr_iu_csr_mtval_30_) );
	DFFPOSX1 DFFPOSX1_1453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_6722__31_), .Q(csr_gpr_iu_csr_mtval_31_) );
	DFFPOSX1 DFFPOSX1_1454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_6710__0_), .Q(csr_gpr_iu_csr_mideleg_0_) );
	DFFPOSX1 DFFPOSX1_1455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_6710__1_), .Q(csr_gpr_iu_csr_mideleg_1_) );
	DFFPOSX1 DFFPOSX1_1456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_6710__2_), .Q(csr_gpr_iu_csr_mideleg_2_) );
	DFFPOSX1 DFFPOSX1_1457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_6710__3_), .Q(csr_gpr_iu_csr_mideleg_3_) );
	DFFPOSX1 DFFPOSX1_1458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_6710__4_), .Q(csr_gpr_iu_csr_mideleg_4_) );
	DFFPOSX1 DFFPOSX1_1459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_6710__5_), .Q(csr_gpr_iu_csr_mideleg_5_) );
	DFFPOSX1 DFFPOSX1_1460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_6710__6_), .Q(csr_gpr_iu_csr_mideleg_6_) );
	DFFPOSX1 DFFPOSX1_1461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_6710__7_), .Q(csr_gpr_iu_csr_mideleg_7_) );
	DFFPOSX1 DFFPOSX1_1462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_6710__8_), .Q(csr_gpr_iu_csr_mideleg_8_) );
	DFFPOSX1 DFFPOSX1_1463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_6710__9_), .Q(csr_gpr_iu_csr_mideleg_9_) );
	DFFPOSX1 DFFPOSX1_1464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_6710__10_), .Q(csr_gpr_iu_csr_mideleg_10_) );
	DFFPOSX1 DFFPOSX1_1465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_6710__11_), .Q(csr_gpr_iu_csr_mideleg_11_) );
	DFFPOSX1 DFFPOSX1_1466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_6710__12_), .Q(csr_gpr_iu_csr_mideleg_12_) );
	DFFPOSX1 DFFPOSX1_1467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_6710__13_), .Q(csr_gpr_iu_csr_mideleg_13_) );
	DFFPOSX1 DFFPOSX1_1468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_6710__14_), .Q(csr_gpr_iu_csr_mideleg_14_) );
	DFFPOSX1 DFFPOSX1_1469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_6710__15_), .Q(csr_gpr_iu_csr_mideleg_15_) );
	DFFPOSX1 DFFPOSX1_1470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_6710__16_), .Q(csr_gpr_iu_csr_mideleg_16_) );
	DFFPOSX1 DFFPOSX1_1471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_6710__17_), .Q(csr_gpr_iu_csr_mideleg_17_) );
	DFFPOSX1 DFFPOSX1_1472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_6710__18_), .Q(csr_gpr_iu_csr_mideleg_18_) );
	DFFPOSX1 DFFPOSX1_1473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_6710__19_), .Q(csr_gpr_iu_csr_mideleg_19_) );
	DFFPOSX1 DFFPOSX1_1474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_6710__20_), .Q(csr_gpr_iu_csr_mideleg_20_) );
	DFFPOSX1 DFFPOSX1_1475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_6710__21_), .Q(csr_gpr_iu_csr_mideleg_21_) );
	DFFPOSX1 DFFPOSX1_1476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_6710__22_), .Q(csr_gpr_iu_csr_mideleg_22_) );
	DFFPOSX1 DFFPOSX1_1477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_6710__23_), .Q(csr_gpr_iu_csr_mideleg_23_) );
	DFFPOSX1 DFFPOSX1_1478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_6710__24_), .Q(csr_gpr_iu_csr_mideleg_24_) );
	DFFPOSX1 DFFPOSX1_1479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_6710__25_), .Q(csr_gpr_iu_csr_mideleg_25_) );
	DFFPOSX1 DFFPOSX1_1480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_6710__26_), .Q(csr_gpr_iu_csr_mideleg_26_) );
	DFFPOSX1 DFFPOSX1_1481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_6710__27_), .Q(csr_gpr_iu_csr_mideleg_27_) );
	DFFPOSX1 DFFPOSX1_1482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_6710__28_), .Q(csr_gpr_iu_csr_mideleg_28_) );
	DFFPOSX1 DFFPOSX1_1483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_6710__29_), .Q(csr_gpr_iu_csr_mideleg_29_) );
	DFFPOSX1 DFFPOSX1_1484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_6710__30_), .Q(csr_gpr_iu_csr_mideleg_30_) );
	DFFPOSX1 DFFPOSX1_1485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_6710__31_), .Q(csr_gpr_iu_csr_mideleg_31_) );
	DFFPOSX1 DFFPOSX1_1486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_6706__0_), .Q(csr_gpr_iu_csr_medeleg_0_) );
	DFFPOSX1 DFFPOSX1_1487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_6706__1_), .Q(csr_gpr_iu_csr_medeleg_1_) );
	DFFPOSX1 DFFPOSX1_1488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_6706__2_), .Q(csr_gpr_iu_csr_medeleg_2_) );
	DFFPOSX1 DFFPOSX1_1489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_6706__3_), .Q(csr_gpr_iu_csr_medeleg_3_) );
	DFFPOSX1 DFFPOSX1_1490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_6706__4_), .Q(csr_gpr_iu_csr_medeleg_4_) );
	DFFPOSX1 DFFPOSX1_1491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_6706__5_), .Q(csr_gpr_iu_csr_medeleg_5_) );
	DFFPOSX1 DFFPOSX1_1492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_6706__6_), .Q(csr_gpr_iu_csr_medeleg_6_) );
	DFFPOSX1 DFFPOSX1_1493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_6706__7_), .Q(csr_gpr_iu_csr_medeleg_7_) );
	DFFPOSX1 DFFPOSX1_1494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_6706__8_), .Q(csr_gpr_iu_csr_medeleg_8_) );
	DFFPOSX1 DFFPOSX1_1495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_6706__9_), .Q(csr_gpr_iu_csr_medeleg_9_) );
	DFFPOSX1 DFFPOSX1_1496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_6706__10_), .Q(csr_gpr_iu_csr_medeleg_10_) );
	DFFPOSX1 DFFPOSX1_1497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_6706__11_), .Q(csr_gpr_iu_csr_medeleg_11_) );
	DFFPOSX1 DFFPOSX1_1498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_6706__12_), .Q(csr_gpr_iu_csr_medeleg_12_) );
	DFFPOSX1 DFFPOSX1_1499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_6706__13_), .Q(csr_gpr_iu_csr_medeleg_13_) );
	DFFPOSX1 DFFPOSX1_1500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6706__14_), .Q(csr_gpr_iu_csr_medeleg_14_) );
	DFFPOSX1 DFFPOSX1_1501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6706__15_), .Q(csr_gpr_iu_csr_medeleg_15_) );
	DFFPOSX1 DFFPOSX1_1502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6706__16_), .Q(csr_gpr_iu_csr_medeleg_16_) );
	DFFPOSX1 DFFPOSX1_1503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6706__17_), .Q(csr_gpr_iu_csr_medeleg_17_) );
	DFFPOSX1 DFFPOSX1_1504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6706__18_), .Q(csr_gpr_iu_csr_medeleg_18_) );
	DFFPOSX1 DFFPOSX1_1505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6706__19_), .Q(csr_gpr_iu_csr_medeleg_19_) );
	DFFPOSX1 DFFPOSX1_1506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6706__20_), .Q(csr_gpr_iu_csr_medeleg_20_) );
	DFFPOSX1 DFFPOSX1_1507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6706__21_), .Q(csr_gpr_iu_csr_medeleg_21_) );
	DFFPOSX1 DFFPOSX1_1508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6706__22_), .Q(csr_gpr_iu_csr_medeleg_22_) );
	DFFPOSX1 DFFPOSX1_1509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6706__23_), .Q(csr_gpr_iu_csr_medeleg_23_) );
	DFFPOSX1 DFFPOSX1_1510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6706__24_), .Q(csr_gpr_iu_csr_medeleg_24_) );
	DFFPOSX1 DFFPOSX1_1511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6706__25_), .Q(csr_gpr_iu_csr_medeleg_25_) );
	DFFPOSX1 DFFPOSX1_1512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6706__26_), .Q(csr_gpr_iu_csr_medeleg_26_) );
	DFFPOSX1 DFFPOSX1_1513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6706__27_), .Q(csr_gpr_iu_csr_medeleg_27_) );
	DFFPOSX1 DFFPOSX1_1514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6706__28_), .Q(csr_gpr_iu_csr_medeleg_28_) );
	DFFPOSX1 DFFPOSX1_1515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_6706__29_), .Q(csr_gpr_iu_csr_medeleg_29_) );
	DFFPOSX1 DFFPOSX1_1516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_6706__30_), .Q(csr_gpr_iu_csr_medeleg_30_) );
	DFFPOSX1 DFFPOSX1_1517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_6706__31_), .Q(csr_gpr_iu_csr_medeleg_31_) );
	DFFPOSX1 DFFPOSX1_1518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_6707_), .Q(csr_gpr_iu_csr_meie) );
	DFFPOSX1 DFFPOSX1_1519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_6740_), .Q(csr_gpr_iu_csr_seie) );
	DFFPOSX1 DFFPOSX1_1520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_6720_), .Q(csr_gpr_iu_csr_mtie) );
	DFFPOSX1 DFFPOSX1_1521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_6749_), .Q(csr_gpr_iu_csr_stie) );
	DFFPOSX1 DFFPOSX1_1522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_6717_), .Q(csr_gpr_iu_csr_msie) );
	DFFPOSX1 DFFPOSX1_1523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_6747_), .Q(csr_gpr_iu_csr_ssie) );
	DFFPOSX1 DFFPOSX1_1524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_6716__0_), .Q(csr_gpr_iu_csr_mscratch_0_) );
	DFFPOSX1 DFFPOSX1_1525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_6716__1_), .Q(csr_gpr_iu_csr_mscratch_1_) );
	DFFPOSX1 DFFPOSX1_1526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_6716__2_), .Q(csr_gpr_iu_csr_mscratch_2_) );
	DFFPOSX1 DFFPOSX1_1527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_6716__3_), .Q(csr_gpr_iu_csr_mscratch_3_) );
	DFFPOSX1 DFFPOSX1_1528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_6716__4_), .Q(csr_gpr_iu_csr_mscratch_4_) );
	DFFPOSX1 DFFPOSX1_1529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_6716__5_), .Q(csr_gpr_iu_csr_mscratch_5_) );
	DFFPOSX1 DFFPOSX1_1530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_6716__6_), .Q(csr_gpr_iu_csr_mscratch_6_) );
	DFFPOSX1 DFFPOSX1_1531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_6716__7_), .Q(csr_gpr_iu_csr_mscratch_7_) );
	DFFPOSX1 DFFPOSX1_1532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_6716__8_), .Q(csr_gpr_iu_csr_mscratch_8_) );
	DFFPOSX1 DFFPOSX1_1533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_6716__9_), .Q(csr_gpr_iu_csr_mscratch_9_) );
	DFFPOSX1 DFFPOSX1_1534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_6716__10_), .Q(csr_gpr_iu_csr_mscratch_10_) );
	DFFPOSX1 DFFPOSX1_1535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_6716__11_), .Q(csr_gpr_iu_csr_mscratch_11_) );
	DFFPOSX1 DFFPOSX1_1536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_6716__12_), .Q(csr_gpr_iu_csr_mscratch_12_) );
	DFFPOSX1 DFFPOSX1_1537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_6716__13_), .Q(csr_gpr_iu_csr_mscratch_13_) );
	DFFPOSX1 DFFPOSX1_1538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_6716__14_), .Q(csr_gpr_iu_csr_mscratch_14_) );
	DFFPOSX1 DFFPOSX1_1539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_6716__15_), .Q(csr_gpr_iu_csr_mscratch_15_) );
	DFFPOSX1 DFFPOSX1_1540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_6716__16_), .Q(csr_gpr_iu_csr_mscratch_16_) );
	DFFPOSX1 DFFPOSX1_1541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_6716__17_), .Q(csr_gpr_iu_csr_mscratch_17_) );
	DFFPOSX1 DFFPOSX1_1542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_6716__18_), .Q(csr_gpr_iu_csr_mscratch_18_) );
	DFFPOSX1 DFFPOSX1_1543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6716__19_), .Q(csr_gpr_iu_csr_mscratch_19_) );
	DFFPOSX1 DFFPOSX1_1544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6716__20_), .Q(csr_gpr_iu_csr_mscratch_20_) );
	DFFPOSX1 DFFPOSX1_1545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6716__21_), .Q(csr_gpr_iu_csr_mscratch_21_) );
	DFFPOSX1 DFFPOSX1_1546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6716__22_), .Q(csr_gpr_iu_csr_mscratch_22_) );
	DFFPOSX1 DFFPOSX1_1547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6716__23_), .Q(csr_gpr_iu_csr_mscratch_23_) );
	DFFPOSX1 DFFPOSX1_1548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6716__24_), .Q(csr_gpr_iu_csr_mscratch_24_) );
	DFFPOSX1 DFFPOSX1_1549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6716__25_), .Q(csr_gpr_iu_csr_mscratch_25_) );
	DFFPOSX1 DFFPOSX1_1550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6716__26_), .Q(csr_gpr_iu_csr_mscratch_26_) );
	DFFPOSX1 DFFPOSX1_1551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6716__27_), .Q(csr_gpr_iu_csr_mscratch_27_) );
	DFFPOSX1 DFFPOSX1_1552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6716__28_), .Q(csr_gpr_iu_csr_mscratch_28_) );
	DFFPOSX1 DFFPOSX1_1553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6716__29_), .Q(csr_gpr_iu_csr_mscratch_29_) );
	DFFPOSX1 DFFPOSX1_1554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6716__30_), .Q(csr_gpr_iu_csr_mscratch_30_) );
	DFFPOSX1 DFFPOSX1_1555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6716__31_), .Q(csr_gpr_iu_csr_mscratch_31_) );
	DFFPOSX1 DFFPOSX1_1556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6726__0_), .Q(csr_gpr_iu_csr_pmp0cfg_0_) );
	DFFPOSX1 DFFPOSX1_1557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6726__1_), .Q(csr_gpr_iu_csr_pmp0cfg_1_) );
	DFFPOSX1 DFFPOSX1_1558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6726__2_), .Q(csr_gpr_iu_csr_pmp0cfg_2_) );
	DFFPOSX1 DFFPOSX1_1559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6726__3_), .Q(csr_gpr_iu_csr_pmp0cfg_3_) );
	DFFPOSX1 DFFPOSX1_1560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6726__4_), .Q(csr_gpr_iu_csr_pmp0cfg_4_) );
	DFFPOSX1 DFFPOSX1_1561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6726__5_), .Q(csr_gpr_iu_csr_pmp0cfg_5_) );
	DFFPOSX1 DFFPOSX1_1562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6726__6_), .Q(csr_gpr_iu_csr_pmp0cfg_6_) );
	DFFPOSX1 DFFPOSX1_1563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6726__7_), .Q(csr_gpr_iu_csr_pmp0cfg_7_) );
	DFFPOSX1 DFFPOSX1_1564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6727__0_), .Q(csr_gpr_iu_csr_pmp1cfg_0_) );
	DFFPOSX1 DFFPOSX1_1565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6727__1_), .Q(csr_gpr_iu_csr_pmp1cfg_1_) );
	DFFPOSX1 DFFPOSX1_1566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6727__2_), .Q(csr_gpr_iu_csr_pmp1cfg_2_) );
	DFFPOSX1 DFFPOSX1_1567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6727__3_), .Q(csr_gpr_iu_csr_pmp1cfg_3_) );
	DFFPOSX1 DFFPOSX1_1568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6727__4_), .Q(csr_gpr_iu_csr_pmp1cfg_4_) );
	DFFPOSX1 DFFPOSX1_1569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6727__5_), .Q(csr_gpr_iu_csr_pmp1cfg_5_) );
	DFFPOSX1 DFFPOSX1_1570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6727__6_), .Q(csr_gpr_iu_csr_pmp1cfg_6_) );
	DFFPOSX1 DFFPOSX1_1571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6727__7_), .Q(csr_gpr_iu_csr_pmp1cfg_7_) );
	DFFPOSX1 DFFPOSX1_1572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6728__0_), .Q(csr_gpr_iu_csr_pmp2cfg_0_) );
	DFFPOSX1 DFFPOSX1_1573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6728__1_), .Q(csr_gpr_iu_csr_pmp2cfg_1_) );
	DFFPOSX1 DFFPOSX1_1574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6728__2_), .Q(csr_gpr_iu_csr_pmp2cfg_2_) );
	DFFPOSX1 DFFPOSX1_1575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6728__3_), .Q(csr_gpr_iu_csr_pmp2cfg_3_) );
	DFFPOSX1 DFFPOSX1_1576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_6728__4_), .Q(csr_gpr_iu_csr_pmp2cfg_4_) );
	DFFPOSX1 DFFPOSX1_1577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_6728__5_), .Q(csr_gpr_iu_csr_pmp2cfg_5_) );
	DFFPOSX1 DFFPOSX1_1578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_6728__6_), .Q(csr_gpr_iu_csr_pmp2cfg_6_) );
	DFFPOSX1 DFFPOSX1_1579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_6728__7_), .Q(csr_gpr_iu_csr_pmp2cfg_7_) );
	DFFPOSX1 DFFPOSX1_1580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_6729__0_), .Q(csr_gpr_iu_csr_pmp3cfg_0_) );
	DFFPOSX1 DFFPOSX1_1581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_6729__1_), .Q(csr_gpr_iu_csr_pmp3cfg_1_) );
	DFFPOSX1 DFFPOSX1_1582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_6729__2_), .Q(csr_gpr_iu_csr_pmp3cfg_2_) );
	DFFPOSX1 DFFPOSX1_1583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_6729__3_), .Q(csr_gpr_iu_csr_pmp3cfg_3_) );
	DFFPOSX1 DFFPOSX1_1584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_6729__4_), .Q(csr_gpr_iu_csr_pmp3cfg_4_) );
	DFFPOSX1 DFFPOSX1_1585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_6729__5_), .Q(csr_gpr_iu_csr_pmp3cfg_5_) );
	DFFPOSX1 DFFPOSX1_1586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_6729__6_), .Q(csr_gpr_iu_csr_pmp3cfg_6_) );
	DFFPOSX1 DFFPOSX1_1587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_6729__7_), .Q(csr_gpr_iu_csr_pmp3cfg_7_) );
	DFFPOSX1 DFFPOSX1_1588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_6730__0_), .Q(csr_gpr_iu_csr_pmp4cfg_0_) );
	DFFPOSX1 DFFPOSX1_1589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_6730__1_), .Q(csr_gpr_iu_csr_pmp4cfg_1_) );
	DFFPOSX1 DFFPOSX1_1590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_6730__2_), .Q(csr_gpr_iu_csr_pmp4cfg_2_) );
	DFFPOSX1 DFFPOSX1_1591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_6730__3_), .Q(csr_gpr_iu_csr_pmp4cfg_3_) );
	DFFPOSX1 DFFPOSX1_1592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6730__4_), .Q(csr_gpr_iu_csr_pmp4cfg_4_) );
	DFFPOSX1 DFFPOSX1_1593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_6730__5_), .Q(csr_gpr_iu_csr_pmp4cfg_5_) );
	DFFPOSX1 DFFPOSX1_1594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_6730__6_), .Q(csr_gpr_iu_csr_pmp4cfg_6_) );
	DFFPOSX1 DFFPOSX1_1595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_6730__7_), .Q(csr_gpr_iu_csr_pmp4cfg_7_) );
	DFFPOSX1 DFFPOSX1_1596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_6731__0_), .Q(csr_gpr_iu_csr_pmp5cfg_0_) );
	DFFPOSX1 DFFPOSX1_1597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_6731__1_), .Q(csr_gpr_iu_csr_pmp5cfg_1_) );
	DFFPOSX1 DFFPOSX1_1598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_6731__2_), .Q(csr_gpr_iu_csr_pmp5cfg_2_) );
	DFFPOSX1 DFFPOSX1_1599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_6731__3_), .Q(csr_gpr_iu_csr_pmp5cfg_3_) );
	DFFPOSX1 DFFPOSX1_1600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6731__4_), .Q(csr_gpr_iu_csr_pmp5cfg_4_) );
	DFFPOSX1 DFFPOSX1_1601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_6731__5_), .Q(csr_gpr_iu_csr_pmp5cfg_5_) );
	DFFPOSX1 DFFPOSX1_1602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_6731__6_), .Q(csr_gpr_iu_csr_pmp5cfg_6_) );
	DFFPOSX1 DFFPOSX1_1603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_6731__7_), .Q(csr_gpr_iu_csr_pmp5cfg_7_) );
	DFFPOSX1 DFFPOSX1_1604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_6732__0_), .Q(csr_gpr_iu_csr_pmp6cfg_0_) );
	DFFPOSX1 DFFPOSX1_1605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_6732__1_), .Q(csr_gpr_iu_csr_pmp6cfg_1_) );
	DFFPOSX1 DFFPOSX1_1606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6732__2_), .Q(csr_gpr_iu_csr_pmp6cfg_2_) );
	DFFPOSX1 DFFPOSX1_1607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6732__3_), .Q(csr_gpr_iu_csr_pmp6cfg_3_) );
	DFFPOSX1 DFFPOSX1_1608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_6732__4_), .Q(csr_gpr_iu_csr_pmp6cfg_4_) );
	DFFPOSX1 DFFPOSX1_1609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6732__5_), .Q(csr_gpr_iu_csr_pmp6cfg_5_) );
	DFFPOSX1 DFFPOSX1_1610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6732__6_), .Q(csr_gpr_iu_csr_pmp6cfg_6_) );
	DFFPOSX1 DFFPOSX1_1611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_6732__7_), .Q(csr_gpr_iu_csr_pmp6cfg_7_) );
	DFFPOSX1 DFFPOSX1_1612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_6733__0_), .Q(csr_gpr_iu_csr_pmp7cfg_0_) );
	DFFPOSX1 DFFPOSX1_1613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_6733__1_), .Q(csr_gpr_iu_csr_pmp7cfg_1_) );
	DFFPOSX1 DFFPOSX1_1614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_6733__2_), .Q(csr_gpr_iu_csr_pmp7cfg_2_) );
	DFFPOSX1 DFFPOSX1_1615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_6733__3_), .Q(csr_gpr_iu_csr_pmp7cfg_3_) );
	DFFPOSX1 DFFPOSX1_1616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_6733__4_), .Q(csr_gpr_iu_csr_pmp7cfg_4_) );
	DFFPOSX1 DFFPOSX1_1617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_6733__5_), .Q(csr_gpr_iu_csr_pmp7cfg_5_) );
	DFFPOSX1 DFFPOSX1_1618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_6733__6_), .Q(csr_gpr_iu_csr_pmp7cfg_6_) );
	DFFPOSX1 DFFPOSX1_1619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_6733__7_), .Q(csr_gpr_iu_csr_pmp7cfg_7_) );
	DFFPOSX1 DFFPOSX1_1620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_6734__0_), .Q(csr_gpr_iu_csr_pmpaddr0_0_) );
	DFFPOSX1 DFFPOSX1_1621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_6734__1_), .Q(csr_gpr_iu_csr_pmpaddr0_1_) );
	DFFPOSX1 DFFPOSX1_1622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_6734__2_), .Q(csr_gpr_iu_csr_pmpaddr0_2_) );
	DFFPOSX1 DFFPOSX1_1623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_6734__3_), .Q(csr_gpr_iu_csr_pmpaddr0_3_) );
	DFFPOSX1 DFFPOSX1_1624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_6734__4_), .Q(csr_gpr_iu_csr_pmpaddr0_4_) );
	DFFPOSX1 DFFPOSX1_1625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_6734__5_), .Q(csr_gpr_iu_csr_pmpaddr0_5_) );
	DFFPOSX1 DFFPOSX1_1626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_6734__6_), .Q(csr_gpr_iu_csr_pmpaddr0_6_) );
	DFFPOSX1 DFFPOSX1_1627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_6734__7_), .Q(csr_gpr_iu_csr_pmpaddr0_7_) );
	DFFPOSX1 DFFPOSX1_1628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_6734__8_), .Q(csr_gpr_iu_csr_pmpaddr0_8_) );
	DFFPOSX1 DFFPOSX1_1629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_6734__9_), .Q(csr_gpr_iu_csr_pmpaddr0_9_) );
	DFFPOSX1 DFFPOSX1_1630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_6734__10_), .Q(csr_gpr_iu_csr_pmpaddr0_10_) );
	DFFPOSX1 DFFPOSX1_1631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_6734__11_), .Q(csr_gpr_iu_csr_pmpaddr0_11_) );
	DFFPOSX1 DFFPOSX1_1632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_6734__12_), .Q(csr_gpr_iu_csr_pmpaddr0_12_) );
	DFFPOSX1 DFFPOSX1_1633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_6734__13_), .Q(csr_gpr_iu_csr_pmpaddr0_13_) );
	DFFPOSX1 DFFPOSX1_1634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_6734__14_), .Q(csr_gpr_iu_csr_pmpaddr0_14_) );
	DFFPOSX1 DFFPOSX1_1635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_6734__15_), .Q(csr_gpr_iu_csr_pmpaddr0_15_) );
	DFFPOSX1 DFFPOSX1_1636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_6734__16_), .Q(csr_gpr_iu_csr_pmpaddr0_16_) );
	DFFPOSX1 DFFPOSX1_1637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_6734__17_), .Q(csr_gpr_iu_csr_pmpaddr0_17_) );
	DFFPOSX1 DFFPOSX1_1638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_6734__18_), .Q(csr_gpr_iu_csr_pmpaddr0_18_) );
	DFFPOSX1 DFFPOSX1_1639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_6734__19_), .Q(csr_gpr_iu_csr_pmpaddr0_19_) );
	DFFPOSX1 DFFPOSX1_1640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_6734__20_), .Q(csr_gpr_iu_csr_pmpaddr0_20_) );
	DFFPOSX1 DFFPOSX1_1641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_6734__21_), .Q(csr_gpr_iu_csr_pmpaddr0_21_) );
	DFFPOSX1 DFFPOSX1_1642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_6734__22_), .Q(csr_gpr_iu_csr_pmpaddr0_22_) );
	DFFPOSX1 DFFPOSX1_1643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_6734__23_), .Q(csr_gpr_iu_csr_pmpaddr0_23_) );
	DFFPOSX1 DFFPOSX1_1644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_6734__24_), .Q(csr_gpr_iu_csr_pmpaddr0_24_) );
	DFFPOSX1 DFFPOSX1_1645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_6734__25_), .Q(csr_gpr_iu_csr_pmpaddr0_25_) );
	DFFPOSX1 DFFPOSX1_1646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_6734__26_), .Q(csr_gpr_iu_csr_pmpaddr0_26_) );
	DFFPOSX1 DFFPOSX1_1647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_6734__27_), .Q(csr_gpr_iu_csr_pmpaddr0_27_) );
	DFFPOSX1 DFFPOSX1_1648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_6734__28_), .Q(csr_gpr_iu_csr_pmpaddr0_28_) );
	DFFPOSX1 DFFPOSX1_1649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_6734__29_), .Q(csr_gpr_iu_csr_pmpaddr0_29_) );
	DFFPOSX1 DFFPOSX1_1650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_6734__30_), .Q(csr_gpr_iu_csr_pmpaddr0_30_) );
	DFFPOSX1 DFFPOSX1_1651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_6734__31_), .Q(csr_gpr_iu_csr_pmpaddr0_31_) );
	DFFPOSX1 DFFPOSX1_1652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_6735__0_), .Q(csr_gpr_iu_csr_pmpaddr1_0_) );
	DFFPOSX1 DFFPOSX1_1653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_6735__1_), .Q(csr_gpr_iu_csr_pmpaddr1_1_) );
	DFFPOSX1 DFFPOSX1_1654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_6735__2_), .Q(csr_gpr_iu_csr_pmpaddr1_2_) );
	DFFPOSX1 DFFPOSX1_1655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_6735__3_), .Q(csr_gpr_iu_csr_pmpaddr1_3_) );
	DFFPOSX1 DFFPOSX1_1656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_6735__4_), .Q(csr_gpr_iu_csr_pmpaddr1_4_) );
	DFFPOSX1 DFFPOSX1_1657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_6735__5_), .Q(csr_gpr_iu_csr_pmpaddr1_5_) );
	DFFPOSX1 DFFPOSX1_1658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_6735__6_), .Q(csr_gpr_iu_csr_pmpaddr1_6_) );
	DFFPOSX1 DFFPOSX1_1659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_6735__7_), .Q(csr_gpr_iu_csr_pmpaddr1_7_) );
	DFFPOSX1 DFFPOSX1_1660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_6735__8_), .Q(csr_gpr_iu_csr_pmpaddr1_8_) );
	DFFPOSX1 DFFPOSX1_1661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6735__9_), .Q(csr_gpr_iu_csr_pmpaddr1_9_) );
	DFFPOSX1 DFFPOSX1_1662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6735__10_), .Q(csr_gpr_iu_csr_pmpaddr1_10_) );
	DFFPOSX1 DFFPOSX1_1663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6735__11_), .Q(csr_gpr_iu_csr_pmpaddr1_11_) );
	DFFPOSX1 DFFPOSX1_1664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6735__12_), .Q(csr_gpr_iu_csr_pmpaddr1_12_) );
	DFFPOSX1 DFFPOSX1_1665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6735__13_), .Q(csr_gpr_iu_csr_pmpaddr1_13_) );
	DFFPOSX1 DFFPOSX1_1666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6735__14_), .Q(csr_gpr_iu_csr_pmpaddr1_14_) );
	DFFPOSX1 DFFPOSX1_1667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6735__15_), .Q(csr_gpr_iu_csr_pmpaddr1_15_) );
	DFFPOSX1 DFFPOSX1_1668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6735__16_), .Q(csr_gpr_iu_csr_pmpaddr1_16_) );
	DFFPOSX1 DFFPOSX1_1669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6735__17_), .Q(csr_gpr_iu_csr_pmpaddr1_17_) );
	DFFPOSX1 DFFPOSX1_1670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6735__18_), .Q(csr_gpr_iu_csr_pmpaddr1_18_) );
	DFFPOSX1 DFFPOSX1_1671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6735__19_), .Q(csr_gpr_iu_csr_pmpaddr1_19_) );
	DFFPOSX1 DFFPOSX1_1672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6735__20_), .Q(csr_gpr_iu_csr_pmpaddr1_20_) );
	DFFPOSX1 DFFPOSX1_1673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6735__21_), .Q(csr_gpr_iu_csr_pmpaddr1_21_) );
	DFFPOSX1 DFFPOSX1_1674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6735__22_), .Q(csr_gpr_iu_csr_pmpaddr1_22_) );
	DFFPOSX1 DFFPOSX1_1675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6735__23_), .Q(csr_gpr_iu_csr_pmpaddr1_23_) );
	DFFPOSX1 DFFPOSX1_1676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_6735__24_), .Q(csr_gpr_iu_csr_pmpaddr1_24_) );
	DFFPOSX1 DFFPOSX1_1677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_6735__25_), .Q(csr_gpr_iu_csr_pmpaddr1_25_) );
	DFFPOSX1 DFFPOSX1_1678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_6735__26_), .Q(csr_gpr_iu_csr_pmpaddr1_26_) );
	DFFPOSX1 DFFPOSX1_1679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_6735__27_), .Q(csr_gpr_iu_csr_pmpaddr1_27_) );
	DFFPOSX1 DFFPOSX1_1680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_6735__28_), .Q(csr_gpr_iu_csr_pmpaddr1_28_) );
	DFFPOSX1 DFFPOSX1_1681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_6735__29_), .Q(csr_gpr_iu_csr_pmpaddr1_29_) );
	DFFPOSX1 DFFPOSX1_1682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_6735__30_), .Q(csr_gpr_iu_csr_pmpaddr1_30_) );
	DFFPOSX1 DFFPOSX1_1683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_6735__31_), .Q(csr_gpr_iu_csr_pmpaddr1_31_) );
	DFFPOSX1 DFFPOSX1_1684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_6736__0_), .Q(csr_gpr_iu_csr_pmpaddr2_0_) );
	DFFPOSX1 DFFPOSX1_1685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_6736__1_), .Q(csr_gpr_iu_csr_pmpaddr2_1_) );
	DFFPOSX1 DFFPOSX1_1686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_6736__2_), .Q(csr_gpr_iu_csr_pmpaddr2_2_) );
	DFFPOSX1 DFFPOSX1_1687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_6736__3_), .Q(csr_gpr_iu_csr_pmpaddr2_3_) );
	DFFPOSX1 DFFPOSX1_1688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_6736__4_), .Q(csr_gpr_iu_csr_pmpaddr2_4_) );
	DFFPOSX1 DFFPOSX1_1689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_6736__5_), .Q(csr_gpr_iu_csr_pmpaddr2_5_) );
	DFFPOSX1 DFFPOSX1_1690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_6736__6_), .Q(csr_gpr_iu_csr_pmpaddr2_6_) );
	DFFPOSX1 DFFPOSX1_1691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_6736__7_), .Q(csr_gpr_iu_csr_pmpaddr2_7_) );
	DFFPOSX1 DFFPOSX1_1692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_6736__8_), .Q(csr_gpr_iu_csr_pmpaddr2_8_) );
	DFFPOSX1 DFFPOSX1_1693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_6736__9_), .Q(csr_gpr_iu_csr_pmpaddr2_9_) );
	DFFPOSX1 DFFPOSX1_1694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_6736__10_), .Q(csr_gpr_iu_csr_pmpaddr2_10_) );
	DFFPOSX1 DFFPOSX1_1695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_6736__11_), .Q(csr_gpr_iu_csr_pmpaddr2_11_) );
	DFFPOSX1 DFFPOSX1_1696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_6736__12_), .Q(csr_gpr_iu_csr_pmpaddr2_12_) );
	DFFPOSX1 DFFPOSX1_1697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_6736__13_), .Q(csr_gpr_iu_csr_pmpaddr2_13_) );
	DFFPOSX1 DFFPOSX1_1698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_6736__14_), .Q(csr_gpr_iu_csr_pmpaddr2_14_) );
	DFFPOSX1 DFFPOSX1_1699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_6736__15_), .Q(csr_gpr_iu_csr_pmpaddr2_15_) );
	DFFPOSX1 DFFPOSX1_1700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_6736__16_), .Q(csr_gpr_iu_csr_pmpaddr2_16_) );
	DFFPOSX1 DFFPOSX1_1701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_6736__17_), .Q(csr_gpr_iu_csr_pmpaddr2_17_) );
	DFFPOSX1 DFFPOSX1_1702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_6736__18_), .Q(csr_gpr_iu_csr_pmpaddr2_18_) );
	DFFPOSX1 DFFPOSX1_1703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_6736__19_), .Q(csr_gpr_iu_csr_pmpaddr2_19_) );
	DFFPOSX1 DFFPOSX1_1704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6736__20_), .Q(csr_gpr_iu_csr_pmpaddr2_20_) );
	DFFPOSX1 DFFPOSX1_1705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6736__21_), .Q(csr_gpr_iu_csr_pmpaddr2_21_) );
	DFFPOSX1 DFFPOSX1_1706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6736__22_), .Q(csr_gpr_iu_csr_pmpaddr2_22_) );
	DFFPOSX1 DFFPOSX1_1707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6736__23_), .Q(csr_gpr_iu_csr_pmpaddr2_23_) );
	DFFPOSX1 DFFPOSX1_1708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6736__24_), .Q(csr_gpr_iu_csr_pmpaddr2_24_) );
	DFFPOSX1 DFFPOSX1_1709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6736__25_), .Q(csr_gpr_iu_csr_pmpaddr2_25_) );
	DFFPOSX1 DFFPOSX1_1710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6736__26_), .Q(csr_gpr_iu_csr_pmpaddr2_26_) );
	DFFPOSX1 DFFPOSX1_1711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6736__27_), .Q(csr_gpr_iu_csr_pmpaddr2_27_) );
	DFFPOSX1 DFFPOSX1_1712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6736__28_), .Q(csr_gpr_iu_csr_pmpaddr2_28_) );
	DFFPOSX1 DFFPOSX1_1713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6736__29_), .Q(csr_gpr_iu_csr_pmpaddr2_29_) );
	DFFPOSX1 DFFPOSX1_1714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6736__30_), .Q(csr_gpr_iu_csr_pmpaddr2_30_) );
	DFFPOSX1 DFFPOSX1_1715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6736__31_), .Q(csr_gpr_iu_csr_pmpaddr2_31_) );
	DFFPOSX1 DFFPOSX1_1716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6737__0_), .Q(csr_gpr_iu_csr_pmpaddr3_0_) );
	DFFPOSX1 DFFPOSX1_1717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6737__1_), .Q(csr_gpr_iu_csr_pmpaddr3_1_) );
	DFFPOSX1 DFFPOSX1_1718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6737__2_), .Q(csr_gpr_iu_csr_pmpaddr3_2_) );
	DFFPOSX1 DFFPOSX1_1719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6737__3_), .Q(csr_gpr_iu_csr_pmpaddr3_3_) );
	DFFPOSX1 DFFPOSX1_1720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6737__4_), .Q(csr_gpr_iu_csr_pmpaddr3_4_) );
	DFFPOSX1 DFFPOSX1_1721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6737__5_), .Q(csr_gpr_iu_csr_pmpaddr3_5_) );
	DFFPOSX1 DFFPOSX1_1722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6737__6_), .Q(csr_gpr_iu_csr_pmpaddr3_6_) );
	DFFPOSX1 DFFPOSX1_1723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6737__7_), .Q(csr_gpr_iu_csr_pmpaddr3_7_) );
	DFFPOSX1 DFFPOSX1_1724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6737__8_), .Q(csr_gpr_iu_csr_pmpaddr3_8_) );
	DFFPOSX1 DFFPOSX1_1725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6737__9_), .Q(csr_gpr_iu_csr_pmpaddr3_9_) );
	DFFPOSX1 DFFPOSX1_1726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6737__10_), .Q(csr_gpr_iu_csr_pmpaddr3_10_) );
	DFFPOSX1 DFFPOSX1_1727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6737__11_), .Q(csr_gpr_iu_csr_pmpaddr3_11_) );
	DFFPOSX1 DFFPOSX1_1728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6737__12_), .Q(csr_gpr_iu_csr_pmpaddr3_12_) );
	DFFPOSX1 DFFPOSX1_1729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6737__13_), .Q(csr_gpr_iu_csr_pmpaddr3_13_) );
	DFFPOSX1 DFFPOSX1_1730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6737__14_), .Q(csr_gpr_iu_csr_pmpaddr3_14_) );
	DFFPOSX1 DFFPOSX1_1731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6737__15_), .Q(csr_gpr_iu_csr_pmpaddr3_15_) );
	DFFPOSX1 DFFPOSX1_1732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6737__16_), .Q(csr_gpr_iu_csr_pmpaddr3_16_) );
	DFFPOSX1 DFFPOSX1_1733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6737__17_), .Q(csr_gpr_iu_csr_pmpaddr3_17_) );
	DFFPOSX1 DFFPOSX1_1734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6737__18_), .Q(csr_gpr_iu_csr_pmpaddr3_18_) );
	DFFPOSX1 DFFPOSX1_1735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6737__19_), .Q(csr_gpr_iu_csr_pmpaddr3_19_) );
	DFFPOSX1 DFFPOSX1_1736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6737__20_), .Q(csr_gpr_iu_csr_pmpaddr3_20_) );
	DFFPOSX1 DFFPOSX1_1737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_6737__21_), .Q(csr_gpr_iu_csr_pmpaddr3_21_) );
	DFFPOSX1 DFFPOSX1_1738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_6737__22_), .Q(csr_gpr_iu_csr_pmpaddr3_22_) );
	DFFPOSX1 DFFPOSX1_1739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_6737__23_), .Q(csr_gpr_iu_csr_pmpaddr3_23_) );
	DFFPOSX1 DFFPOSX1_1740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_6737__24_), .Q(csr_gpr_iu_csr_pmpaddr3_24_) );
	DFFPOSX1 DFFPOSX1_1741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_6737__25_), .Q(csr_gpr_iu_csr_pmpaddr3_25_) );
	DFFPOSX1 DFFPOSX1_1742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_6737__26_), .Q(csr_gpr_iu_csr_pmpaddr3_26_) );
	DFFPOSX1 DFFPOSX1_1743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_6737__27_), .Q(csr_gpr_iu_csr_pmpaddr3_27_) );
	DFFPOSX1 DFFPOSX1_1744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_6737__28_), .Q(csr_gpr_iu_csr_pmpaddr3_28_) );
	DFFPOSX1 DFFPOSX1_1745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_6737__29_), .Q(csr_gpr_iu_csr_pmpaddr3_29_) );
	DFFPOSX1 DFFPOSX1_1746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_6737__30_), .Q(csr_gpr_iu_csr_pmpaddr3_30_) );
	DFFPOSX1 DFFPOSX1_1747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_6737__31_), .Q(csr_gpr_iu_csr_pmpaddr3_31_) );
	DFFPOSX1 DFFPOSX1_1748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_6752__0_), .Q(csr_gpr_iu_csr_stvec_0_) );
	DFFPOSX1 DFFPOSX1_1749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_6752__1_), .Q(csr_gpr_iu_csr_stvec_1_) );
	DFFPOSX1 DFFPOSX1_1750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_6752__2_), .Q(csr_gpr_iu_csr_stvec_2_) );
	DFFPOSX1 DFFPOSX1_1751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_6752__3_), .Q(csr_gpr_iu_csr_stvec_3_) );
	DFFPOSX1 DFFPOSX1_1752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_6752__4_), .Q(csr_gpr_iu_csr_stvec_4_) );
	DFFPOSX1 DFFPOSX1_1753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_6752__5_), .Q(csr_gpr_iu_csr_stvec_5_) );
	DFFPOSX1 DFFPOSX1_1754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_6752__6_), .Q(csr_gpr_iu_csr_stvec_6_) );
	DFFPOSX1 DFFPOSX1_1755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_6752__7_), .Q(csr_gpr_iu_csr_stvec_7_) );
	DFFPOSX1 DFFPOSX1_1756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_6752__8_), .Q(csr_gpr_iu_csr_stvec_8_) );
	DFFPOSX1 DFFPOSX1_1757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_6752__9_), .Q(csr_gpr_iu_csr_stvec_9_) );
	DFFPOSX1 DFFPOSX1_1758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_6752__10_), .Q(csr_gpr_iu_csr_stvec_10_) );
	DFFPOSX1 DFFPOSX1_1759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_6752__11_), .Q(csr_gpr_iu_csr_stvec_11_) );
	DFFPOSX1 DFFPOSX1_1760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_6752__12_), .Q(csr_gpr_iu_csr_stvec_12_) );
	DFFPOSX1 DFFPOSX1_1761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6752__13_), .Q(csr_gpr_iu_csr_stvec_13_) );
	DFFPOSX1 DFFPOSX1_1762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_6752__14_), .Q(csr_gpr_iu_csr_stvec_14_) );
	DFFPOSX1 DFFPOSX1_1763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_6752__15_), .Q(csr_gpr_iu_csr_stvec_15_) );
	DFFPOSX1 DFFPOSX1_1764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_6752__16_), .Q(csr_gpr_iu_csr_stvec_16_) );
	DFFPOSX1 DFFPOSX1_1765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_6752__17_), .Q(csr_gpr_iu_csr_stvec_17_) );
	DFFPOSX1 DFFPOSX1_1766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_6752__18_), .Q(csr_gpr_iu_csr_stvec_18_) );
	DFFPOSX1 DFFPOSX1_1767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6752__19_), .Q(csr_gpr_iu_csr_stvec_19_) );
	DFFPOSX1 DFFPOSX1_1768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6752__20_), .Q(csr_gpr_iu_csr_stvec_20_) );
	DFFPOSX1 DFFPOSX1_1769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_6752__21_), .Q(csr_gpr_iu_csr_stvec_21_) );
	DFFPOSX1 DFFPOSX1_1770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6752__22_), .Q(csr_gpr_iu_csr_stvec_22_) );
	DFFPOSX1 DFFPOSX1_1771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_6752__23_), .Q(csr_gpr_iu_csr_stvec_23_) );
	DFFPOSX1 DFFPOSX1_1772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_6752__24_), .Q(csr_gpr_iu_csr_stvec_24_) );
	DFFPOSX1 DFFPOSX1_1773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_6752__25_), .Q(csr_gpr_iu_csr_stvec_25_) );
	DFFPOSX1 DFFPOSX1_1774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_6752__26_), .Q(csr_gpr_iu_csr_stvec_26_) );
	DFFPOSX1 DFFPOSX1_1775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_6752__27_), .Q(csr_gpr_iu_csr_stvec_27_) );
	DFFPOSX1 DFFPOSX1_1776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_6752__28_), .Q(csr_gpr_iu_csr_stvec_28_) );
	DFFPOSX1 DFFPOSX1_1777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_6752__29_), .Q(csr_gpr_iu_csr_stvec_29_) );
	DFFPOSX1 DFFPOSX1_1778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_6752__30_), .Q(csr_gpr_iu_csr_stvec_30_) );
	DFFPOSX1 DFFPOSX1_1779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_6752__31_), .Q(csr_gpr_iu_csr_stvec_31_) );
	DFFPOSX1 DFFPOSX1_1780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_6751__0_), .Q(csr_gpr_iu_csr_stval_0_) );
	DFFPOSX1 DFFPOSX1_1781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_6751__1_), .Q(csr_gpr_iu_csr_stval_1_) );
	DFFPOSX1 DFFPOSX1_1782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_6751__2_), .Q(csr_gpr_iu_csr_stval_2_) );
	DFFPOSX1 DFFPOSX1_1783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_6751__3_), .Q(csr_gpr_iu_csr_stval_3_) );
	DFFPOSX1 DFFPOSX1_1784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_6751__4_), .Q(csr_gpr_iu_csr_stval_4_) );
	DFFPOSX1 DFFPOSX1_1785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_6751__5_), .Q(csr_gpr_iu_csr_stval_5_) );
	DFFPOSX1 DFFPOSX1_1786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_6751__6_), .Q(csr_gpr_iu_csr_stval_6_) );
	DFFPOSX1 DFFPOSX1_1787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_6751__7_), .Q(csr_gpr_iu_csr_stval_7_) );
	DFFPOSX1 DFFPOSX1_1788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_6751__8_), .Q(csr_gpr_iu_csr_stval_8_) );
	DFFPOSX1 DFFPOSX1_1789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_6751__9_), .Q(csr_gpr_iu_csr_stval_9_) );
	DFFPOSX1 DFFPOSX1_1790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_6751__10_), .Q(csr_gpr_iu_csr_stval_10_) );
	DFFPOSX1 DFFPOSX1_1791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_6751__11_), .Q(csr_gpr_iu_csr_stval_11_) );
	DFFPOSX1 DFFPOSX1_1792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_6751__12_), .Q(csr_gpr_iu_csr_stval_12_) );
	DFFPOSX1 DFFPOSX1_1793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_6751__13_), .Q(csr_gpr_iu_csr_stval_13_) );
	DFFPOSX1 DFFPOSX1_1794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_6751__14_), .Q(csr_gpr_iu_csr_stval_14_) );
	DFFPOSX1 DFFPOSX1_1795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_6751__15_), .Q(csr_gpr_iu_csr_stval_15_) );
	DFFPOSX1 DFFPOSX1_1796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_6751__16_), .Q(csr_gpr_iu_csr_stval_16_) );
	DFFPOSX1 DFFPOSX1_1797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_6751__17_), .Q(csr_gpr_iu_csr_stval_17_) );
	DFFPOSX1 DFFPOSX1_1798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_6751__18_), .Q(csr_gpr_iu_csr_stval_18_) );
	DFFPOSX1 DFFPOSX1_1799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_6751__19_), .Q(csr_gpr_iu_csr_stval_19_) );
	DFFPOSX1 DFFPOSX1_1800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_6751__20_), .Q(csr_gpr_iu_csr_stval_20_) );
	DFFPOSX1 DFFPOSX1_1801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_6751__21_), .Q(csr_gpr_iu_csr_stval_21_) );
	DFFPOSX1 DFFPOSX1_1802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_6751__22_), .Q(csr_gpr_iu_csr_stval_22_) );
	DFFPOSX1 DFFPOSX1_1803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_6751__23_), .Q(csr_gpr_iu_csr_stval_23_) );
	DFFPOSX1 DFFPOSX1_1804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_6751__24_), .Q(csr_gpr_iu_csr_stval_24_) );
	DFFPOSX1 DFFPOSX1_1805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_6751__25_), .Q(csr_gpr_iu_csr_stval_25_) );
	DFFPOSX1 DFFPOSX1_1806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_6751__26_), .Q(csr_gpr_iu_csr_stval_26_) );
	DFFPOSX1 DFFPOSX1_1807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_6751__27_), .Q(csr_gpr_iu_csr_stval_27_) );
	DFFPOSX1 DFFPOSX1_1808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_6751__28_), .Q(csr_gpr_iu_csr_stval_28_) );
	DFFPOSX1 DFFPOSX1_1809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_6751__29_), .Q(csr_gpr_iu_csr_stval_29_) );
	DFFPOSX1 DFFPOSX1_1810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_6751__30_), .Q(csr_gpr_iu_csr_stval_30_) );
	DFFPOSX1 DFFPOSX1_1811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_6751__31_), .Q(csr_gpr_iu_csr_stval_31_) );
	DFFPOSX1 DFFPOSX1_1812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_6742__0_), .Q(csr_gpr_iu_csr_sepc_0_) );
	DFFPOSX1 DFFPOSX1_1813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_6742__1_), .Q(csr_gpr_iu_csr_sepc_1_) );
	DFFPOSX1 DFFPOSX1_1814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_6742__2_), .Q(csr_gpr_iu_csr_sepc_2_) );
	DFFPOSX1 DFFPOSX1_1815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_6742__3_), .Q(csr_gpr_iu_csr_sepc_3_) );
	DFFPOSX1 DFFPOSX1_1816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_6742__4_), .Q(csr_gpr_iu_csr_sepc_4_) );
	DFFPOSX1 DFFPOSX1_1817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_6742__5_), .Q(csr_gpr_iu_csr_sepc_5_) );
	DFFPOSX1 DFFPOSX1_1818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_6742__6_), .Q(csr_gpr_iu_csr_sepc_6_) );
	DFFPOSX1 DFFPOSX1_1819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_6742__7_), .Q(csr_gpr_iu_csr_sepc_7_) );
	DFFPOSX1 DFFPOSX1_1820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_6742__8_), .Q(csr_gpr_iu_csr_sepc_8_) );
	DFFPOSX1 DFFPOSX1_1821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_6742__9_), .Q(csr_gpr_iu_csr_sepc_9_) );
	DFFPOSX1 DFFPOSX1_1822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6742__10_), .Q(csr_gpr_iu_csr_sepc_10_) );
	DFFPOSX1 DFFPOSX1_1823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6742__11_), .Q(csr_gpr_iu_csr_sepc_11_) );
	DFFPOSX1 DFFPOSX1_1824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6742__12_), .Q(csr_gpr_iu_csr_sepc_12_) );
	DFFPOSX1 DFFPOSX1_1825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6742__13_), .Q(csr_gpr_iu_csr_sepc_13_) );
	DFFPOSX1 DFFPOSX1_1826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6742__14_), .Q(csr_gpr_iu_csr_sepc_14_) );
	DFFPOSX1 DFFPOSX1_1827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6742__15_), .Q(csr_gpr_iu_csr_sepc_15_) );
	DFFPOSX1 DFFPOSX1_1828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6742__16_), .Q(csr_gpr_iu_csr_sepc_16_) );
	DFFPOSX1 DFFPOSX1_1829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6742__17_), .Q(csr_gpr_iu_csr_sepc_17_) );
	DFFPOSX1 DFFPOSX1_1830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6742__18_), .Q(csr_gpr_iu_csr_sepc_18_) );
	DFFPOSX1 DFFPOSX1_1831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6742__19_), .Q(csr_gpr_iu_csr_sepc_19_) );
	DFFPOSX1 DFFPOSX1_1832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6742__20_), .Q(csr_gpr_iu_csr_sepc_20_) );
	DFFPOSX1 DFFPOSX1_1833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6742__21_), .Q(csr_gpr_iu_csr_sepc_21_) );
	DFFPOSX1 DFFPOSX1_1834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6742__22_), .Q(csr_gpr_iu_csr_sepc_22_) );
	DFFPOSX1 DFFPOSX1_1835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6742__23_), .Q(csr_gpr_iu_csr_sepc_23_) );
	DFFPOSX1 DFFPOSX1_1836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6742__24_), .Q(csr_gpr_iu_csr_sepc_24_) );
	DFFPOSX1 DFFPOSX1_1837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_6742__25_), .Q(csr_gpr_iu_csr_sepc_25_) );
	DFFPOSX1 DFFPOSX1_1838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_6742__26_), .Q(csr_gpr_iu_csr_sepc_26_) );
	DFFPOSX1 DFFPOSX1_1839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_6742__27_), .Q(csr_gpr_iu_csr_sepc_27_) );
	DFFPOSX1 DFFPOSX1_1840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_6742__28_), .Q(csr_gpr_iu_csr_sepc_28_) );
	DFFPOSX1 DFFPOSX1_1841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_6742__29_), .Q(csr_gpr_iu_csr_sepc_29_) );
	DFFPOSX1 DFFPOSX1_1842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_6742__30_), .Q(csr_gpr_iu_csr_sepc_30_) );
	DFFPOSX1 DFFPOSX1_1843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_6742__31_), .Q(csr_gpr_iu_csr_sepc_31_) );
	DFFPOSX1 DFFPOSX1_1844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_6739__0_), .Q(csr_gpr_iu_csr_scause_0_) );
	DFFPOSX1 DFFPOSX1_1845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_6739__1_), .Q(csr_gpr_iu_csr_scause_1_) );
	DFFPOSX1 DFFPOSX1_1846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_6739__2_), .Q(csr_gpr_iu_csr_scause_2_) );
	DFFPOSX1 DFFPOSX1_1847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_6739__3_), .Q(csr_gpr_iu_csr_scause_3_) );
	DFFPOSX1 DFFPOSX1_1848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_6739__4_), .Q(csr_gpr_iu_csr_scause_4_) );
	DFFPOSX1 DFFPOSX1_1849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_6739__5_), .Q(csr_gpr_iu_csr_scause_5_) );
	DFFPOSX1 DFFPOSX1_1850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_6739__6_), .Q(csr_gpr_iu_csr_scause_6_) );
	DFFPOSX1 DFFPOSX1_1851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_6739__7_), .Q(csr_gpr_iu_csr_scause_7_) );
	DFFPOSX1 DFFPOSX1_1852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_6739__8_), .Q(csr_gpr_iu_csr_scause_8_) );
	DFFPOSX1 DFFPOSX1_1853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_6739__9_), .Q(csr_gpr_iu_csr_scause_9_) );
	DFFPOSX1 DFFPOSX1_1854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_6739__10_), .Q(csr_gpr_iu_csr_scause_10_) );
	DFFPOSX1 DFFPOSX1_1855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_6739__11_), .Q(csr_gpr_iu_csr_scause_11_) );
	DFFPOSX1 DFFPOSX1_1856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_6739__12_), .Q(csr_gpr_iu_csr_scause_12_) );
	DFFPOSX1 DFFPOSX1_1857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_6739__13_), .Q(csr_gpr_iu_csr_scause_13_) );
	DFFPOSX1 DFFPOSX1_1858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_6739__14_), .Q(csr_gpr_iu_csr_scause_14_) );
	DFFPOSX1 DFFPOSX1_1859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_6739__15_), .Q(csr_gpr_iu_csr_scause_15_) );
	DFFPOSX1 DFFPOSX1_1860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_6739__16_), .Q(csr_gpr_iu_csr_scause_16_) );
	DFFPOSX1 DFFPOSX1_1861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_6739__17_), .Q(csr_gpr_iu_csr_scause_17_) );
	DFFPOSX1 DFFPOSX1_1862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_6739__18_), .Q(csr_gpr_iu_csr_scause_18_) );
	DFFPOSX1 DFFPOSX1_1863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_6739__19_), .Q(csr_gpr_iu_csr_scause_19_) );
	DFFPOSX1 DFFPOSX1_1864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_6739__20_), .Q(csr_gpr_iu_csr_scause_20_) );
	DFFPOSX1 DFFPOSX1_1865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6739__21_), .Q(csr_gpr_iu_csr_scause_21_) );
	DFFPOSX1 DFFPOSX1_1866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6739__22_), .Q(csr_gpr_iu_csr_scause_22_) );
	DFFPOSX1 DFFPOSX1_1867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6739__23_), .Q(csr_gpr_iu_csr_scause_23_) );
	DFFPOSX1 DFFPOSX1_1868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6739__24_), .Q(csr_gpr_iu_csr_scause_24_) );
	DFFPOSX1 DFFPOSX1_1869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6739__25_), .Q(csr_gpr_iu_csr_scause_25_) );
	DFFPOSX1 DFFPOSX1_1870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6739__26_), .Q(csr_gpr_iu_csr_scause_26_) );
	DFFPOSX1 DFFPOSX1_1871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6739__27_), .Q(csr_gpr_iu_csr_scause_27_) );
	DFFPOSX1 DFFPOSX1_1872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6739__28_), .Q(csr_gpr_iu_csr_scause_28_) );
	DFFPOSX1 DFFPOSX1_1873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6739__29_), .Q(csr_gpr_iu_csr_scause_29_) );
	DFFPOSX1 DFFPOSX1_1874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6739__30_), .Q(csr_gpr_iu_csr_scause_30_) );
	DFFPOSX1 DFFPOSX1_1875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6739__31_), .Q(csr_gpr_iu_csr_scause_31_) );
	DFFPOSX1 DFFPOSX1_1876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6746__0_), .Q(csr_gpr_iu_csr_sscratch_0_) );
	DFFPOSX1 DFFPOSX1_1877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6746__1_), .Q(csr_gpr_iu_csr_sscratch_1_) );
	DFFPOSX1 DFFPOSX1_1878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6746__2_), .Q(csr_gpr_iu_csr_sscratch_2_) );
	DFFPOSX1 DFFPOSX1_1879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6746__3_), .Q(csr_gpr_iu_csr_sscratch_3_) );
	DFFPOSX1 DFFPOSX1_1880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6746__4_), .Q(csr_gpr_iu_csr_sscratch_4_) );
	DFFPOSX1 DFFPOSX1_1881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6746__5_), .Q(csr_gpr_iu_csr_sscratch_5_) );
	DFFPOSX1 DFFPOSX1_1882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6746__6_), .Q(csr_gpr_iu_csr_sscratch_6_) );
	DFFPOSX1 DFFPOSX1_1883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6746__7_), .Q(csr_gpr_iu_csr_sscratch_7_) );
	DFFPOSX1 DFFPOSX1_1884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6746__8_), .Q(csr_gpr_iu_csr_sscratch_8_) );
	DFFPOSX1 DFFPOSX1_1885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6746__9_), .Q(csr_gpr_iu_csr_sscratch_9_) );
	DFFPOSX1 DFFPOSX1_1886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6746__10_), .Q(csr_gpr_iu_csr_sscratch_10_) );
	DFFPOSX1 DFFPOSX1_1887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6746__11_), .Q(csr_gpr_iu_csr_sscratch_11_) );
	DFFPOSX1 DFFPOSX1_1888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6746__12_), .Q(csr_gpr_iu_csr_sscratch_12_) );
	DFFPOSX1 DFFPOSX1_1889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6746__13_), .Q(csr_gpr_iu_csr_sscratch_13_) );
	DFFPOSX1 DFFPOSX1_1890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6746__14_), .Q(csr_gpr_iu_csr_sscratch_14_) );
	DFFPOSX1 DFFPOSX1_1891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6746__15_), .Q(csr_gpr_iu_csr_sscratch_15_) );
	DFFPOSX1 DFFPOSX1_1892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6746__16_), .Q(csr_gpr_iu_csr_sscratch_16_) );
	DFFPOSX1 DFFPOSX1_1893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6746__17_), .Q(csr_gpr_iu_csr_sscratch_17_) );
	DFFPOSX1 DFFPOSX1_1894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6746__18_), .Q(csr_gpr_iu_csr_sscratch_18_) );
	DFFPOSX1 DFFPOSX1_1895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6746__19_), .Q(csr_gpr_iu_csr_sscratch_19_) );
	DFFPOSX1 DFFPOSX1_1896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6746__20_), .Q(csr_gpr_iu_csr_sscratch_20_) );
	DFFPOSX1 DFFPOSX1_1897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_6746__21_), .Q(csr_gpr_iu_csr_sscratch_21_) );
	DFFPOSX1 DFFPOSX1_1898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_6746__22_), .Q(csr_gpr_iu_csr_sscratch_22_) );
	DFFPOSX1 DFFPOSX1_1899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_6746__23_), .Q(csr_gpr_iu_csr_sscratch_23_) );
	DFFPOSX1 DFFPOSX1_1900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_6746__24_), .Q(csr_gpr_iu_csr_sscratch_24_) );
	DFFPOSX1 DFFPOSX1_1901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_6746__25_), .Q(csr_gpr_iu_csr_sscratch_25_) );
	DFFPOSX1 DFFPOSX1_1902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_6746__26_), .Q(csr_gpr_iu_csr_sscratch_26_) );
	DFFPOSX1 DFFPOSX1_1903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_6746__27_), .Q(csr_gpr_iu_csr_sscratch_27_) );
	DFFPOSX1 DFFPOSX1_1904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_6746__28_), .Q(csr_gpr_iu_csr_sscratch_28_) );
	DFFPOSX1 DFFPOSX1_1905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_6746__29_), .Q(csr_gpr_iu_csr_sscratch_29_) );
	DFFPOSX1 DFFPOSX1_1906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_6746__30_), .Q(csr_gpr_iu_csr_sscratch_30_) );
	DFFPOSX1 DFFPOSX1_1907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_6746__31_), .Q(csr_gpr_iu_csr_sscratch_31_) );
	NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_1_), .B(biu_ins_0_), .Y(_10981_) );
	NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .B(biu_ins_3_), .C(_10981_), .Y(_10982_) );
	NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(biu_ins_6_), .C(biu_ins_5_), .Y(_10819_) );
	NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(_10982_), .Y(_10820_) );
	NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(biu_ins_12_), .Y(_10821_) );
	INVX1 INVX1_1702 ( .gnd(gnd), .vdd(vdd), .A(_10820_), .Y(_10822_) );
	NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10822_), .Y(_10823_) );
	NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(biu_ins_12_), .Y(_10824_) );
	NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(_10824_), .Y(_10825_) );
	INVX1 INVX1_1703 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .Y(_10826_) );
	INVX1 INVX1_1704 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_12_), .Y(_10827_) );
	NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(_10827_), .Y(_10828_) );
	NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_10828_), .B(_10826_), .Y(_10829_) );
	OAI21X1 OAI21X1_4352 ( .gnd(gnd), .vdd(vdd), .A(_10820_), .B(_10829_), .C(_10823_), .Y(biu_exce_chk_opc_2_) );
	INVX1 INVX1_1705 ( .gnd(gnd), .vdd(vdd), .A(_10824_), .Y(_10830_) );
	OAI21X1 OAI21X1_4353 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10824_), .C(_10822_), .Y(_10831_) );
	INVX1 INVX1_1706 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_5_), .Y(_10832_) );
	NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(biu_ins_6_), .C(_10832_), .Y(_10833_) );
	NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10982_), .Y(_10834_) );
	OAI21X1 OAI21X1_4354 ( .gnd(gnd), .vdd(vdd), .A(_10830_), .B(_10834_), .C(_10831_), .Y(biu_exce_chk_opc_0_) );
	INVX1 INVX1_1707 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .Y(_10835_) );
	NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_10835_), .B(_10828_), .Y(_10836_) );
	NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_10820_), .B(_10829_), .Y(_10837_) );
	NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_10830_), .B(_10834_), .Y(_10838_) );
	AOI21X1 AOI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_10838_), .B(biu_ins_13_), .C(_10837_), .Y(_10839_) );
	OAI21X1 OAI21X1_4355 ( .gnd(gnd), .vdd(vdd), .A(_10834_), .B(_10836_), .C(_10839_), .Y(biu_exce_chk_opc_1_) );
	NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(biu_ins_5_), .Y(_10840_) );
	OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_10840_), .B(biu_ins_6_), .Y(_10841_) );
	INVX1 INVX1_1708 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .Y(_10842_) );
	NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_3_), .B(_10842_), .C(_10981_), .Y(_10843_) );
	INVX1 INVX1_1709 ( .gnd(gnd), .vdd(vdd), .A(_10843_), .Y(_10844_) );
	NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_10841_), .B(_10844_), .Y(csr_gpr_iu_ins_dec_lui) );
	INVX1 INVX1_1710 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .Y(_10845_) );
	NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .B(biu_ins_5_), .C(_10845_), .Y(_10846_) );
	INVX1 INVX1_1711 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .Y(_10847_) );
	NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(_10847_), .C(_10832_), .Y(_10848_) );
	NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .B(biu_ins_3_), .Y(_10849_) );
	NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_10981_), .B(_10849_), .Y(_10850_) );
	AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_10848_), .B(_10850_), .Y(csr_gpr_iu_ins_dec_jal) );
	INVX1 INVX1_1712 ( .gnd(gnd), .vdd(vdd), .A(_10848_), .Y(_10851_) );
	NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_10844_), .B(_10851_), .Y(csr_gpr_iu_ins_dec_jalr) );
	NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(_10850_), .Y(_10852_) );
	AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_1_), .B(biu_ins_0_), .Y(_10853_) );
	NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .B(biu_ins_3_), .Y(_10854_) );
	NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_10854_), .B(_10853_), .Y(_10855_) );
	OAI21X1 OAI21X1_4356 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_5_), .B(_10847_), .C(biu_ins_4_), .Y(_10856_) );
	NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_10850_), .B(_10833_), .Y(_10857_) );
	INVX1 INVX1_1713 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .Y(_10858_) );
	NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .B(_10851_), .Y(_10859_) );
	AOI21X1 AOI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_10859_), .B(_10825_), .C(_10858_), .Y(_10860_) );
	OAI21X1 OAI21X1_4357 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .B(_10856_), .C(_10860_), .Y(_10861_) );
	NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(biu_ins_13_), .C(biu_ins_12_), .Y(_10862_) );
	INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .Y(_10863_) );
	AOI22X1 AOI22X1_633 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(_10850_), .C(_10843_), .D(_10848_), .Y(_10864_) );
	OAI21X1 OAI21X1_4358 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(_10833_), .C(_10982_), .Y(_10865_) );
	NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .B(_10845_), .Y(_10866_) );
	AOI22X1 AOI22X1_634 ( .gnd(gnd), .vdd(vdd), .A(_10843_), .B(_10866_), .C(_10848_), .D(_10850_), .Y(_10867_) );
	AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_10867_), .B(_10865_), .Y(_10868_) );
	OAI21X1 OAI21X1_4359 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10864_), .C(_10868_), .Y(_10869_) );
	NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_10869_), .B(_10861_), .Y(csr_gpr_iu_ill_ins) );
	NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .B(_10982_), .C(_10848_), .Y(_10870_) );
	INVX1 INVX1_1714 ( .gnd(gnd), .vdd(vdd), .A(_10870_), .Y(beq) );
	INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(_10859_), .Y(_10871_) );
	NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10871_), .Y(bne) );
	NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(_10821_), .Y(_10872_) );
	NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_10872_), .B(_10871_), .Y(blt) );
	INVX1 INVX1_1715 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .Y(_10873_) );
	NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(biu_ins_12_), .C(_10873_), .Y(_10874_) );
	NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .B(_10871_), .Y(bge) );
	NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(biu_ins_13_), .C(_10827_), .Y(_10875_) );
	NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10871_), .Y(bltu) );
	NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .B(biu_ins_13_), .C(biu_ins_12_), .Y(_10876_) );
	INVX1 INVX1_1716 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .Y(_10877_) );
	NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_10877_), .B(_10982_), .C(_10848_), .Y(_10878_) );
	INVX1 INVX1_1717 ( .gnd(gnd), .vdd(vdd), .A(_10878_), .Y(bgeu) );
	NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf2), .B(biu_ins_29_bF_buf1), .Y(_10879_) );
	NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf3), .B(biu_ins_27_bF_buf2), .Y(_10880_) );
	NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf0), .B(biu_ins_25_bF_buf1), .C(biu_ins_31_bF_buf0), .Y(_10881_) );
	NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(_10879_), .B(_10880_), .C(_10881_), .Y(_10882_) );
	NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(biu_ins_6_), .C(biu_ins_5_), .Y(_10883_) );
	INVX1 INVX1_1718 ( .gnd(gnd), .vdd(vdd), .A(_10883_), .Y(_10884_) );
	NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_10884_), .B(_10982_), .Y(_10885_) );
	OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_10885_), .B(_10863_), .Y(_10886_) );
	NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10886_), .Y(csr_gpr_iu_ecall) );
	INVX1 INVX1_1719 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf0), .Y(_10887_) );
	NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(biu_ins_30_bF_buf1), .C(biu_ins_29_bF_buf0), .Y(_10888_) );
	NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10888_), .Y(_10889_) );
	OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .B(biu_ins_26_bF_buf3), .Y(_10890_) );
	OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_10886_), .B(_10890_), .Y(_10891_) );
	NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_10887_), .B(_10891_), .Y(csr_gpr_iu_ebreak) );
	INVX1 INVX1_1720 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf0), .Y(_10892_) );
	NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .B(_10832_), .Y(_10893_) );
	AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_10982_), .B(_10893_), .Y(_10894_) );
	NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_7_), .B(_10894_), .Y(_10895_) );
	OAI21X1 OAI21X1_4360 ( .gnd(gnd), .vdd(vdd), .A(_10892_), .B(_10894_), .C(_10895_), .Y(csr_gpr_iu_imm12_0_) );
	INVX1 INVX1_1721 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf3), .Y(_10896_) );
	NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .B(_10894_), .Y(_10897_) );
	OAI21X1 OAI21X1_4361 ( .gnd(gnd), .vdd(vdd), .A(_10896_), .B(_10894_), .C(_10897_), .Y(csr_gpr_iu_imm12_1_) );
	INVX1 INVX1_1722 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf1), .Y(_10898_) );
	NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_9_), .B(_10894_), .Y(_10899_) );
	OAI21X1 OAI21X1_4362 ( .gnd(gnd), .vdd(vdd), .A(_10898_), .B(_10894_), .C(_10899_), .Y(csr_gpr_iu_imm12_2_) );
	INVX1 INVX1_1723 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .Y(_10900_) );
	NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_10_), .B(_10894_), .Y(_10901_) );
	OAI21X1 OAI21X1_4363 ( .gnd(gnd), .vdd(vdd), .A(_10900_), .B(_10894_), .C(_10901_), .Y(csr_gpr_iu_imm12_3_) );
	INVX1 INVX1_1724 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_10902_) );
	NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .B(_10894_), .Y(_10903_) );
	OAI21X1 OAI21X1_4364 ( .gnd(gnd), .vdd(vdd), .A(_10902_), .B(_10894_), .C(_10903_), .Y(csr_gpr_iu_imm12_4_) );
	NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .B(_10840_), .Y(_10904_) );
	NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(_10853_), .B(_10854_), .C(_10904_), .Y(_10905_) );
	NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10905_), .Y(csr_gpr_iu_ins_dec_sllp) );
	NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .B(_10905_), .Y(csr_gpr_iu_ins_dec_sltp) );
	NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(biu_ins_12_), .C(_10835_), .Y(_10906_) );
	NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_10906_), .B(_10905_), .Y(csr_gpr_iu_ins_dec_sltup) );
	NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_10872_), .B(_10905_), .Y(csr_gpr_iu_ins_dec_xorp) );
	NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_10846_), .B(_10982_), .Y(_10907_) );
	NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10907_), .Y(csr_gpr_iu_ins_dec_ori) );
	NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .B(_10907_), .Y(andi) );
	NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10907_), .Y(csr_gpr_iu_ins_dec_slli) );
	NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_10906_), .B(_10885_), .Y(csr_gpr_iu_csrrc) );
	NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .B(_10885_), .Y(csr_gpr_iu_csrrwi) );
	NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10885_), .Y(csr_gpr_iu_csrrsi) );
	NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .B(_10885_), .Y(csr_gpr_iu_csrrci) );
	NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10905_), .Y(csr_gpr_iu_ins_dec_orp) );
	NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .B(_10905_), .Y(andp) );
	NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10885_), .Y(csr_gpr_iu_csrrw) );
	NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .B(_10885_), .Y(csr_gpr_iu_csrrs) );
	INVX1 INVX1_1725 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .Y(_10908_) );
	NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(_10846_), .B(_10982_), .C(_10908_), .Y(_10909_) );
	NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10909_), .Y(csr_gpr_iu_ins_dec_srli) );
	INVX1 INVX1_1726 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf0), .Y(_10910_) );
	NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf3), .B(_10910_), .Y(_10911_) );
	NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10881_), .C(_10911_), .Y(_10912_) );
	NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10909_), .Y(csr_gpr_iu_ins_dec_srai) );
	NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10907_), .Y(addi) );
	NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .B(_10907_), .Y(csr_gpr_iu_ins_dec_slti) );
	NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_10906_), .B(_10907_), .Y(csr_gpr_iu_ins_dec_sltiu) );
	NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .B(_10855_), .C(_10841_), .Y(_10913_) );
	NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10905_), .Y(_10914_) );
	NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10912_), .Y(_10915_) );
	OAI21X1 OAI21X1_4365 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10914_), .C(_10915_), .Y(_10916_) );
	AOI21X1 AOI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10876_), .C(_10905_), .Y(_10917_) );
	AOI21X1 AOI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10836_), .C(_10907_), .Y(_10918_) );
	NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_10917_), .B(_10918_), .Y(_10919_) );
	AOI21X1 AOI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .B(_10906_), .C(_10907_), .Y(_10920_) );
	AOI21X1 AOI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(biu_ins_12_), .C(_10824_), .Y(_10921_) );
	NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(_10921_), .B(_10982_), .C(_10848_), .Y(_10922_) );
	OAI21X1 OAI21X1_4366 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10885_), .C(_10922_), .Y(_10923_) );
	NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_10920_), .B(_10923_), .Y(_10924_) );
	NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_10916_), .B(_10919_), .C(_10924_), .Y(_10925_) );
	NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(_10870_), .B(_10864_), .C(_10867_), .Y(_10926_) );
	AOI21X1 AOI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10912_), .C(_10909_), .Y(_10927_) );
	NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_10927_), .B(_10926_), .Y(_10928_) );
	AOI21X1 AOI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_10907_), .B(_10905_), .C(_10872_), .Y(_10929_) );
	AOI21X1 AOI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_10876_), .C(_10907_), .Y(_10930_) );
	NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_10930_), .B(_10929_), .Y(_10931_) );
	OAI21X1 OAI21X1_4367 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10905_), .C(_10878_), .Y(_10932_) );
	AOI21X1 AOI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_10825_), .B(_10906_), .C(_10905_), .Y(_10933_) );
	NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_10933_), .B(_10932_), .Y(_10934_) );
	NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_10931_), .B(_10934_), .C(_10928_), .Y(_10935_) );
	NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .B(_10935_), .Y(csr_gpr_iu_ins_dec_ins_flow_0_) );
	INVX1 INVX1_1727 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf1), .Y(_10936_) );
	NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(_10936_), .Y(_10937_) );
	NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf2), .B(_10879_), .C(_10937_), .Y(_10938_) );
	NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_10938_), .B(_10857_), .Y(csr_gpr_iu_ins_dec_sc_w) );
	NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(_10857_), .Y(_10939_) );
	INVX1 INVX1_1728 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf1), .Y(_10940_) );
	NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf0), .B(_10940_), .Y(_10941_) );
	AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_10941_), .B(_10879_), .Y(_10942_) );
	AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .B(_10942_), .Y(csr_gpr_iu_ins_dec_lr_w) );
	OAI21X1 OAI21X1_4368 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .B(_10938_), .C(_10865_), .Y(_10943_) );
	AOI21X1 AOI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .B(_10942_), .C(_10943_), .Y(csr_gpr_iu_ins_dec_ins_flow_1_) );
	NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_10879_), .B(_10880_), .Y(_10944_) );
	NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(_10858_), .Y(_10945_) );
	NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_10944_), .B(_10945_), .Y(amomin) );
	INVX1 INVX1_1729 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf2), .Y(_10946_) );
	NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf3), .B(_10946_), .Y(_10947_) );
	NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10947_), .Y(_10948_) );
	NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_10948_), .B(_10945_), .Y(amomax) );
	AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_10911_), .B(_10880_), .Y(_10949_) );
	INVX1 INVX1_1730 ( .gnd(gnd), .vdd(vdd), .A(_10949_), .Y(_10950_) );
	NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_10950_), .B(_10945_), .Y(amominu) );
	NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_10910_), .B(_10946_), .Y(_10951_) );
	NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10951_), .Y(_10952_) );
	NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10945_), .Y(amomaxu) );
	INVX1 INVX1_1731 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .Y(_10953_) );
	NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_10948_), .B(_10953_), .Y(amoxor) );
	NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_10940_), .B(_10879_), .C(_10937_), .Y(_10954_) );
	NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_10954_), .B(_10857_), .Y(amoswap) );
	NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .B(_10857_), .Y(amoadd) );
	NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10953_), .Y(amoand) );
	INVX1 INVX1_1732 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf2), .Y(_10955_) );
	NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(_10955_), .B(_10880_), .C(_10951_), .Y(_10956_) );
	AOI21X1 AOI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_10956_), .B(_10889_), .C(_10857_), .Y(_10957_) );
	NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(_10955_), .B(_10880_), .C(_10947_), .Y(_10958_) );
	AOI21X1 AOI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_10954_), .B(_10958_), .C(_10857_), .Y(_10959_) );
	NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_10959_), .B(_10957_), .Y(_10960_) );
	NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(_10880_), .C(_10911_), .Y(_10961_) );
	NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(_10880_), .C(_10951_), .Y(_10962_) );
	AOI21X1 AOI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_10962_), .B(_10961_), .C(_10857_), .Y(_10963_) );
	NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(_10879_), .C(_10880_), .Y(_10964_) );
	NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(_10880_), .C(_10947_), .Y(_10965_) );
	AOI21X1 AOI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_10965_), .B(_10964_), .C(_10857_), .Y(_10966_) );
	NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_10966_), .B(_10963_), .Y(_10967_) );
	NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(_10967_), .B(_10960_), .C(csr_gpr_iu_ins_dec_ins_flow_1_), .Y(_10968_) );
	NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .B(_10968_), .C(_10935_), .Y(csr_gpr_iu_ins_dec_ins_flow_3_) );
	INVX1 INVX1_1733 ( .gnd(gnd), .vdd(vdd), .A(_10914_), .Y(_10969_) );
	NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10969_), .Y(addp) );
	NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10969_), .Y(csr_gpr_iu_ins_dec_subp) );
	INVX1 INVX1_1734 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .Y(_10970_) );
	NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10970_), .Y(csr_gpr_iu_ins_dec_srlp) );
	NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10970_), .Y(csr_gpr_iu_ins_dec_srap) );
	NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_10950_), .B(_10953_), .Y(amoor) );
	INVX1 INVX1_1735 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .Y(_10971_) );
	NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf2), .B(_10887_), .C(_10971_), .Y(_10972_) );
	NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_10972_), .B(_10886_), .Y(csr_gpr_iu_csr_ret) );
	NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10820_), .Y(csr_gpr_iu_ins_dec_lb) );
	NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10820_), .Y(csr_gpr_iu_ins_dec_lh) );
	NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10885_), .Y(csr_gpr_iu_csr_csr_wr) );
	NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(_10838_), .Y(_10973_) );
	NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(biu_exce_chk_statu_cpu_2_), .Y(_10974_) );
	AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(biu_exce_chk_statu_cpu_0_), .Y(_10975_) );
	NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_10974_), .B(_10975_), .C(_10852_), .Y(_10976_) );
	NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .B(_10835_), .Y(_10977_) );
	AOI21X1 AOI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_10859_), .B(_10977_), .C(_10976_), .Y(_10978_) );
	NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(_10973_), .B(_10978_), .C(_10891_), .Y(_10979_) );
	AOI21X1 AOI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_10830_), .B(_10836_), .C(_10834_), .Y(_10980_) );
	AOI21X1 AOI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_10839_), .B(_10980_), .C(_10979_), .Y(csr_gpr_iu_gpr_wr) );
	INVX1 INVX1_1736 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .Y(_10986_) );
	NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(_10986_), .Y(_10987_) );
	INVX1 INVX1_1737 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .Y(_10988_) );
	NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(_10988_), .Y(_10989_) );
	AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10989_), .Y(csr_gpr_iu_csr_meip_wr) );
	INVX1 INVX1_1738 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_4_), .Y(_10990_) );
	NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf2), .B(biu_mmu_msu_1_), .Y(_10991_) );
	NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_timer_int), .B(_10991_), .Y(_10992_) );
	INVX1 INVX1_1739 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_timer_int), .Y(_10993_) );
	INVX1 INVX1_1740 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_sti), .Y(_10994_) );
	NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf2), .B(biu_ins_20_bF_buf6), .Y(_10995_) );
	NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf3), .B(biu_ins_25_bF_buf3), .Y(_10996_) );
	AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_10995_), .B(_10996_), .Y(_10997_) );
	AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf1), .B(biu_mmu_msu_1_), .Y(_10998_) );
	NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .B(biu_ins_23_), .Y(_10999_) );
	NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .B(_10999_), .C(_10997_), .Y(_11000_) );
	INVX1 INVX1_1741 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf0), .Y(_11001_) );
	NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(_11001_), .Y(_11002_) );
	NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf2), .B(biu_ins_29_bF_buf1), .Y(_11003_) );
	NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf0), .B(biu_ins_26_bF_buf1), .C(csr_gpr_iu_csr_csr_wr), .Y(_11004_) );
	INVX1 INVX1_1742 ( .gnd(gnd), .vdd(vdd), .A(_11004_), .Y(_11005_) );
	NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_11003_), .B(_11002_), .C(_11005_), .Y(_11006_) );
	NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .B(_11000_), .Y(_11007_) );
	MUX2X1 MUX2X1_166 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(csr_gpr_iu_csr_stip), .S(_11007_), .Y(_11008_) );
	NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .B(_10994_), .C(_11008_), .Y(_11009_) );
	INVX1 INVX1_1743 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf0), .Y(_11010_) );
	NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .B(_11010_), .Y(_11011_) );
	NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_sie), .B(_11011_), .Y(_11012_) );
	NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_stie), .B(csr_gpr_iu_csr_mideleg_5_), .Y(_11013_) );
	NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_11013_), .B(_11012_), .Y(_11014_) );
	NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_11014_), .B(_11009_), .Y(_11015_) );
	OAI21X1 OAI21X1_4369 ( .gnd(gnd), .vdd(vdd), .A(_10990_), .B(_10992_), .C(_11015_), .Y(csr_gpr_iu_int_ctrl_sti) );
	NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .B(_11008_), .Y(csr_gpr_iu_csr_stip_in) );
	INVX1 INVX1_1744 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_ext_int), .Y(_11016_) );
	INVX1 INVX1_1745 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .Y(_11017_) );
	NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seip), .B(_11007_), .Y(_11018_) );
	AOI21X1 AOI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_11017_), .B(_11007_), .C(_11018_), .Y(_11019_) );
	NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_sei), .B(_11019_), .Y(_11020_) );
	NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_8_), .B(csr_gpr_iu_int_ctrl_ext_int), .C(_10991_), .Y(_11021_) );
	INVX1 INVX1_1746 ( .gnd(gnd), .vdd(vdd), .A(_11012_), .Y(_11022_) );
	NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_seie), .B(csr_gpr_iu_csr_mideleg_9_), .C(_11022_), .Y(_11023_) );
	AOI22X1 AOI22X1_635 ( .gnd(gnd), .vdd(vdd), .A(_11021_), .B(_11023_), .C(_11016_), .D(_11020_), .Y(csr_gpr_iu_int_ctrl_sei) );
	INVX1 INVX1_1747 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .Y(csr_gpr_iu_csr_seip_in) );
	INVX1 INVX1_1748 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_soft_int), .Y(_11024_) );
	INVX1 INVX1_1749 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_ssi), .Y(_11025_) );
	MUX2X1 MUX2X1_167 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(csr_gpr_iu_csr_ssip), .S(_11007_), .Y(_11026_) );
	NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(_11024_), .B(_11025_), .C(_11026_), .Y(_11027_) );
	INVX1 INVX1_1750 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_0_), .Y(_11028_) );
	NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_soft_int), .B(_10991_), .Y(_11029_) );
	NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_ssie), .B(csr_gpr_iu_csr_mideleg_1_), .C(_11022_), .Y(_11030_) );
	OAI21X1 OAI21X1_4370 ( .gnd(gnd), .vdd(vdd), .A(_11028_), .B(_11029_), .C(_11030_), .Y(_11031_) );
	AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_11027_), .B(_11031_), .Y(csr_gpr_iu_int_ctrl_ssi) );
	NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_11025_), .B(_11026_), .Y(csr_gpr_iu_csr_ssip_in) );
	INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_1_), .Y(_11032_) );
	INVX1 INVX1_1751 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_9_), .Y(_11033_) );
	NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf4), .B(_11032_), .C(_11033_), .Y(_11034_) );
	INVX1 INVX1_1752 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_8_), .Y(_11035_) );
	NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_11035_), .B(_10991_), .Y(_11036_) );
	AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mie), .B(csr_gpr_iu_csr_meie), .Y(_11037_) );
	NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .B(_11037_), .Y(_11038_) );
	NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(_11034_), .B(_11036_), .C(_11038_), .Y(_11039_) );
	NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_ext_int), .B(_11039_), .Y(_11040_) );
	INVX1 INVX1_1753 ( .gnd(gnd), .vdd(vdd), .A(_11040_), .Y(csr_gpr_iu_csr_meip_in) );
	INVX1 INVX1_1754 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_2_), .Y(_11041_) );
	INVX1 INVX1_1755 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_5_), .Y(_11042_) );
	AOI22X1 AOI22X1_636 ( .gnd(gnd), .vdd(vdd), .A(_11041_), .B(csr_gpr_iu_ill_ins), .C(csr_gpr_iu_int_ctrl_load_acc_fault), .D(_11042_), .Y(_11043_) );
	INVX1 INVX1_1756 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_4_), .Y(_11044_) );
	INVX1 INVX1_1757 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_6_), .Y(_11045_) );
	AOI22X1 AOI22X1_637 ( .gnd(gnd), .vdd(vdd), .A(_11044_), .B(csr_gpr_iu_int_ctrl_load_addr_mis), .C(csr_gpr_iu_int_ctrl_st_addr_mis), .D(_11045_), .Y(_11046_) );
	INVX1 INVX1_1758 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_0_), .Y(_11047_) );
	INVX1 INVX1_1759 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_1_), .Y(_11048_) );
	AOI22X1 AOI22X1_638 ( .gnd(gnd), .vdd(vdd), .A(_11047_), .B(csr_gpr_iu_ins_addr_mis), .C(csr_gpr_iu_ins_acc_fault), .D(_11048_), .Y(_11049_) );
	NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11046_), .C(_11049_), .Y(_11050_) );
	INVX1 INVX1_1760 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_page_fault), .Y(_11051_) );
	INVX1 INVX1_1761 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_ld_page_fault), .Y(_11052_) );
	OAI22X1 OAI22X1_814 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_13_), .B(_11052_), .C(_11051_), .D(csr_gpr_iu_csr_medeleg_15_), .Y(_11053_) );
	INVX1 INVX1_1762 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .Y(_11054_) );
	INVX1 INVX1_1763 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_acc_fault), .Y(_11055_) );
	OAI22X1 OAI22X1_815 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_7_), .B(_11055_), .C(_11054_), .D(csr_gpr_iu_csr_medeleg_12_), .Y(_11056_) );
	OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_11053_), .B(_11056_), .Y(_11057_) );
	NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_11050_), .B(_11057_), .Y(_11058_) );
	INVX1 INVX1_1764 ( .gnd(gnd), .vdd(vdd), .A(_11058_), .Y(_11059_) );
	INVX4 INVX4_32 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ecall), .Y(_11060_) );
	INVX1 INVX1_1765 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ebreak), .Y(_11061_) );
	OAI22X1 OAI22X1_816 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_3_), .B(_11061_), .C(csr_gpr_iu_csr_medeleg_8_), .D(_11060_), .Y(_11062_) );
	OAI21X1 OAI21X1_4371 ( .gnd(gnd), .vdd(vdd), .A(_11062_), .B(_11059_), .C(_10991_), .Y(_11063_) );
	NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ecall), .B(_10998_), .Y(_11064_) );
	INVX1 INVX1_1766 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_addr_mis), .Y(_11065_) );
	NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_acc_fault), .B(csr_gpr_iu_ins_addr_mis), .Y(_11066_) );
	NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_11065_), .B(_11066_), .Y(_11067_) );
	NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(csr_gpr_iu_int_ctrl_st_acc_fault), .Y(_11068_) );
	OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_load_acc_fault), .B(csr_gpr_iu_int_ctrl_load_addr_mis), .Y(_11069_) );
	INVX1 INVX1_1767 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .Y(_11070_) );
	NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_page_fault), .B(csr_gpr_iu_int_ctrl_ld_page_fault), .Y(_11071_) );
	NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ill_ins), .B(csr_gpr_iu_ebreak), .Y(_11072_) );
	AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_11071_), .B(_11072_), .Y(_11073_) );
	NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(_11068_), .B(_11070_), .C(_11073_), .Y(_11074_) );
	OAI21X1 OAI21X1_4372 ( .gnd(gnd), .vdd(vdd), .A(_11067_), .B(_11074_), .C(_10998_), .Y(_11075_) );
	NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_11064_), .B(_11075_), .Y(_11076_) );
	INVX1 INVX1_1768 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_3_), .Y(_11077_) );
	INVX1 INVX1_1769 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_9_), .Y(_11078_) );
	AOI22X1 AOI22X1_639 ( .gnd(gnd), .vdd(vdd), .A(_11077_), .B(csr_gpr_iu_ebreak), .C(csr_gpr_iu_ecall), .D(_11078_), .Y(_11079_) );
	NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_11079_), .B(_11058_), .Y(_11080_) );
	AOI21X1 AOI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_11080_), .B(_11011_), .C(_11076_), .Y(_11081_) );
	AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_11081_), .B(_11063_), .Y(_11082_) );
	AOI22X1 AOI22X1_640 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_page_fault), .B(csr_gpr_iu_csr_medeleg_15_), .C(csr_gpr_iu_int_ctrl_ld_page_fault), .D(csr_gpr_iu_csr_medeleg_13_), .Y(_11083_) );
	AOI22X1 AOI22X1_641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_load_acc_fault), .B(csr_gpr_iu_csr_medeleg_5_), .C(csr_gpr_iu_ill_ins), .D(csr_gpr_iu_csr_medeleg_2_), .Y(_11084_) );
	AOI22X1 AOI22X1_642 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_addr_mis), .B(csr_gpr_iu_csr_medeleg_6_), .C(csr_gpr_iu_int_ctrl_load_addr_mis), .D(csr_gpr_iu_csr_medeleg_4_), .Y(_11085_) );
	AOI22X1 AOI22X1_643 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_acc_fault), .B(csr_gpr_iu_csr_medeleg_1_), .C(csr_gpr_iu_ins_addr_mis), .D(csr_gpr_iu_csr_medeleg_0_), .Y(_11086_) );
	NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_11085_), .C(_11086_), .Y(_11087_) );
	INVX1 INVX1_1770 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .Y(_11088_) );
	AOI22X1 AOI22X1_644 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(csr_gpr_iu_csr_medeleg_12_), .C(csr_gpr_iu_int_ctrl_st_acc_fault), .D(csr_gpr_iu_csr_medeleg_7_), .Y(_11089_) );
	NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_11083_), .B(_11089_), .C(_11088_), .Y(_11090_) );
	INVX1 INVX1_1771 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_8_), .Y(_11091_) );
	NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_medeleg_3_), .B(csr_gpr_iu_ebreak), .Y(_11092_) );
	OAI21X1 OAI21X1_4373 ( .gnd(gnd), .vdd(vdd), .A(_11091_), .B(_11060_), .C(_11092_), .Y(_11093_) );
	OAI21X1 OAI21X1_4374 ( .gnd(gnd), .vdd(vdd), .A(_11093_), .B(_11090_), .C(_10991_), .Y(_11094_) );
	OAI21X1 OAI21X1_4375 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11078_), .C(_11092_), .Y(_11095_) );
	OAI21X1 OAI21X1_4376 ( .gnd(gnd), .vdd(vdd), .A(_11095_), .B(_11090_), .C(_11011_), .Y(_11096_) );
	NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_11094_), .B(_11096_), .Y(_11097_) );
	INVX1 INVX1_1772 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_1_), .Y(_11098_) );
	NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf3), .B(_11032_), .C(_11098_), .Y(_11099_) );
	NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_11028_), .B(_10991_), .Y(_11100_) );
	NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mie), .B(csr_gpr_iu_csr_msie), .C(_10998_), .Y(_11101_) );
	NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .B(_11100_), .C(_11101_), .Y(_11102_) );
	AOI22X1 AOI22X1_645 ( .gnd(gnd), .vdd(vdd), .A(_11039_), .B(csr_gpr_iu_int_ctrl_ext_int), .C(csr_gpr_iu_int_ctrl_soft_int), .D(_11102_), .Y(_11103_) );
	INVX1 INVX1_1773 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_sei), .Y(_11104_) );
	NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_sti), .B(csr_gpr_iu_int_ctrl_ssi), .Y(_11105_) );
	NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_11104_), .B(_11105_), .Y(_11106_) );
	NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_10990_), .B(_10991_), .Y(_11107_) );
	AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mie), .B(csr_gpr_iu_csr_mtie), .Y(_11108_) );
	NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .B(_11108_), .Y(_11109_) );
	INVX1 INVX1_1774 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_mideleg_5_), .Y(_11110_) );
	NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf2), .B(_11032_), .C(_11110_), .Y(_11111_) );
	NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_11111_), .B(_11107_), .C(_11109_), .Y(_11112_) );
	NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_timer_int), .B(_11112_), .Y(_11113_) );
	INVX1 INVX1_1775 ( .gnd(gnd), .vdd(vdd), .A(_11113_), .Y(csr_gpr_iu_csr_mtip_in) );
	NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_11106_), .B(csr_gpr_iu_csr_mtip_in), .Y(_11114_) );
	NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_11103_), .B(_11114_), .Y(csr_gpr_iu_int_acc) );
	NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .B(csr_gpr_iu_int_acc), .Y(_11115_) );
	NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_11115_), .B(_11082_), .Y(csr_gpr_iu_csr_priv_d_0_) );
	AOI22X1 AOI22X1_646 ( .gnd(gnd), .vdd(vdd), .A(_11104_), .B(_11105_), .C(csr_gpr_iu_int_ctrl_timer_int), .D(_11112_), .Y(_11116_) );
	AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_11103_), .B(_11116_), .Y(_11117_) );
	OAI21X1 OAI21X1_4377 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .B(_11117_), .C(_11082_), .Y(csr_gpr_iu_csr_priv_d_1_) );
	NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_soft_int), .B(_11102_), .Y(_11118_) );
	INVX1 INVX1_1776 ( .gnd(gnd), .vdd(vdd), .A(_11118_), .Y(csr_gpr_iu_csr_msip_in) );
	INVX8 INVX8_90 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ill_ins), .Y(_11119_) );
	INVX1 INVX1_1777 ( .gnd(gnd), .vdd(vdd), .A(_10991_), .Y(_11120_) );
	NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11120_), .Y(_11121_) );
	AOI21X1 AOI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf1), .B(csr_gpr_iu_ecall), .C(csr_gpr_iu_int_ctrl_st_acc_fault), .Y(_11122_) );
	OAI21X1 OAI21X1_4378 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11121_), .C(_11122_), .Y(_11123_) );
	AOI21X1 AOI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .B(_11065_), .C(csr_gpr_iu_int_ctrl_load_acc_fault), .Y(_11124_) );
	OAI21X1 OAI21X1_4379 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_load_addr_mis), .B(_11124_), .C(_11061_), .Y(_11125_) );
	AOI21X1 AOI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_11125_), .B(_11119__bF_buf4), .C(csr_gpr_iu_ins_acc_fault), .Y(_11126_) );
	NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_addr_mis), .B(_11126_), .Y(csr_gpr_iu_cause_0_) );
	INVX8 INVX8_91 ( .gnd(gnd), .vdd(vdd), .A(_11066_), .Y(_11127_) );
	NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_11051_), .B(_11116_), .C(_11103_), .Y(_11128_) );
	NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(csr_gpr_iu_int_ctrl_ld_page_fault), .Y(_11129_) );
	INVX1 INVX1_1778 ( .gnd(gnd), .vdd(vdd), .A(_11129_), .Y(_11130_) );
	NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ecall), .B(_11011_), .Y(_11131_) );
	OAI21X1 OAI21X1_4380 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11120_), .C(_11131_), .Y(_11132_) );
	NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_11130_), .B(_11132_), .Y(_11133_) );
	AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_11128_), .B(_11133_), .Y(_11134_) );
	NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_11055_), .B(_11065_), .C(_11064_), .Y(_11135_) );
	OAI21X1 OAI21X1_4381 ( .gnd(gnd), .vdd(vdd), .A(_11135_), .B(_11134_), .C(_11070_), .Y(_11136_) );
	AOI21X1 AOI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_11136_), .B(_11072_), .C(_11127__bF_buf4), .Y(csr_gpr_iu_cause_1_) );
	NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_11066_), .B(_11072_), .Y(_11137_) );
	OAI21X1 OAI21X1_4382 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_sei), .B(csr_gpr_iu_int_ctrl_ssi), .C(_10994_), .Y(_11138_) );
	AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_11103_), .B(_11138_), .Y(_11139_) );
	NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_int_ctrl_st_page_fault), .B(csr_gpr_iu_csr_mtip_in), .Y(_11140_) );
	NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_11129_), .B(_11140_), .Y(_11141_) );
	INVX1 INVX1_1779 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .Y(_11142_) );
	NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_11142_), .B(_11121_), .Y(_11143_) );
	OAI21X1 OAI21X1_4383 ( .gnd(gnd), .vdd(vdd), .A(_11139_), .B(_11141_), .C(_11143_), .Y(_11144_) );
	NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_11055_), .B(_11065_), .Y(_11145_) );
	NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_11145_), .Y(_11146_) );
	AOI21X1 AOI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_11144_), .B(_11146_), .C(_11137_), .Y(csr_gpr_iu_cause_2_) );
	AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11118_), .Y(_11147_) );
	OAI21X1 OAI21X1_4384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_meip_in), .B(_11105_), .C(_11147_), .Y(_11148_) );
	OAI21X1 OAI21X1_4385 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11120_), .C(_11054_), .Y(_11149_) );
	OAI21X1 OAI21X1_4386 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .B(_11060_), .C(_11071_), .Y(_11150_) );
	NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_11150_), .B(_11149_), .Y(_11151_) );
	NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(_11066_), .B(_11072_), .C(_11146_), .Y(_11152_) );
	AOI21X1 AOI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_11148_), .B(_11151_), .C(_11152_), .Y(csr_gpr_iu_cause_3_) );
	NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_11067_), .B(_11074_), .Y(_11153_) );
	OAI21X1 OAI21X1_4387 ( .gnd(gnd), .vdd(vdd), .A(biu_mmu_msu_0_bF_buf0), .B(_11032_), .C(csr_gpr_iu_ecall), .Y(_11154_) );
	NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_11154_), .B(_11153_), .Y(_11155_) );
	INVX1 INVX1_1780 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .Y(csr_gpr_iu_cause_27_) );
	NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(csr_gpr_iu_int_acc), .Y(csr_gpr_iu_cause_31_) );
	NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .B(_11066_), .Y(_11156_) );
	NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_11071_), .B(_11146_), .Y(_11157_) );
	INVX8 INVX8_92 ( .gnd(gnd), .vdd(vdd), .A(_11157_), .Y(_11158_) );
	INVX1 INVX1_1781 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_0_), .Y(_11159_) );
	OAI21X1 OAI21X1_4388 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11159_), .C(_11158__bF_buf7), .Y(_11160_) );
	OAI21X1 OAI21X1_4389 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_11158__bF_buf6), .C(_11160_), .Y(_11161_) );
	OAI21X1 OAI21X1_4390 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf3), .C(biu_pc_0_), .Y(_11162_) );
	OAI21X1 OAI21X1_4391 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11161_), .C(_11162_), .Y(csr_gpr_iu_csr_tval_0_) );
	INVX1 INVX1_1782 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_1_), .Y(_11163_) );
	OAI21X1 OAI21X1_4392 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11163_), .C(_11158__bF_buf5), .Y(_11164_) );
	OAI21X1 OAI21X1_4393 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_11158__bF_buf4), .C(_11164_), .Y(_11165_) );
	OAI21X1 OAI21X1_4394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf2), .C(biu_pc_1_), .Y(_11166_) );
	OAI21X1 OAI21X1_4395 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11165_), .C(_11166_), .Y(csr_gpr_iu_csr_tval_1_) );
	INVX1 INVX1_1783 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_2_), .Y(_11167_) );
	OAI21X1 OAI21X1_4396 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11167_), .C(_11158__bF_buf3), .Y(_11168_) );
	OAI21X1 OAI21X1_4397 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_2_), .B(_11158__bF_buf2), .C(_11168_), .Y(_11169_) );
	OAI21X1 OAI21X1_4398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(_11127__bF_buf1), .C(biu_pc_2_), .Y(_11170_) );
	OAI21X1 OAI21X1_4399 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11169_), .C(_11170_), .Y(csr_gpr_iu_csr_tval_2_) );
	INVX1 INVX1_1784 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_3_), .Y(_11171_) );
	OAI21X1 OAI21X1_4400 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11171_), .C(_11158__bF_buf1), .Y(_11172_) );
	OAI21X1 OAI21X1_4401 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_3_), .B(_11158__bF_buf0), .C(_11172_), .Y(_11173_) );
	OAI21X1 OAI21X1_4402 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(_11127__bF_buf0), .C(biu_pc_3_), .Y(_11174_) );
	OAI21X1 OAI21X1_4403 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11173_), .C(_11174_), .Y(csr_gpr_iu_csr_tval_3_) );
	INVX1 INVX1_1785 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_4_), .Y(_11175_) );
	OAI21X1 OAI21X1_4404 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11175_), .C(_11158__bF_buf7), .Y(_11176_) );
	OAI21X1 OAI21X1_4405 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_4_), .B(_11158__bF_buf6), .C(_11176_), .Y(_11177_) );
	OAI21X1 OAI21X1_4406 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11127__bF_buf4), .C(biu_pc_4_), .Y(_11178_) );
	OAI21X1 OAI21X1_4407 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11177_), .C(_11178_), .Y(csr_gpr_iu_csr_tval_4_) );
	INVX1 INVX1_1786 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_5_), .Y(_11179_) );
	OAI21X1 OAI21X1_4408 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11179_), .C(_11158__bF_buf5), .Y(_11180_) );
	OAI21X1 OAI21X1_4409 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_5_), .B(_11158__bF_buf4), .C(_11180_), .Y(_11181_) );
	OAI21X1 OAI21X1_4410 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(_11127__bF_buf3), .C(biu_pc_5_), .Y(_11182_) );
	OAI21X1 OAI21X1_4411 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11181_), .C(_11182_), .Y(csr_gpr_iu_csr_tval_5_) );
	INVX1 INVX1_1787 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_6_), .Y(_11183_) );
	OAI21X1 OAI21X1_4412 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11183_), .C(_11158__bF_buf3), .Y(_11184_) );
	OAI21X1 OAI21X1_4413 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_11158__bF_buf2), .C(_11184_), .Y(_11185_) );
	OAI21X1 OAI21X1_4414 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf2), .C(biu_pc_6_), .Y(_11186_) );
	OAI21X1 OAI21X1_4415 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11185_), .C(_11186_), .Y(csr_gpr_iu_csr_tval_6_) );
	INVX1 INVX1_1788 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_7_), .Y(_11187_) );
	OAI21X1 OAI21X1_4416 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11187_), .C(_11158__bF_buf1), .Y(_11188_) );
	OAI21X1 OAI21X1_4417 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_7_), .B(_11158__bF_buf0), .C(_11188_), .Y(_11189_) );
	OAI21X1 OAI21X1_4418 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf1), .C(biu_pc_7_), .Y(_11190_) );
	OAI21X1 OAI21X1_4419 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11189_), .C(_11190_), .Y(csr_gpr_iu_csr_tval_7_) );
	INVX1 INVX1_1789 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_8_), .Y(_11191_) );
	OAI21X1 OAI21X1_4420 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11191_), .C(_11158__bF_buf7), .Y(_11192_) );
	OAI21X1 OAI21X1_4421 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_11158__bF_buf6), .C(_11192_), .Y(_11193_) );
	OAI21X1 OAI21X1_4422 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(_11127__bF_buf0), .C(biu_pc_8_), .Y(_11194_) );
	OAI21X1 OAI21X1_4423 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11193_), .C(_11194_), .Y(csr_gpr_iu_csr_tval_8_) );
	INVX1 INVX1_1790 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_9_), .Y(_11195_) );
	OAI21X1 OAI21X1_4424 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11195_), .C(_11158__bF_buf5), .Y(_11196_) );
	OAI21X1 OAI21X1_4425 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_9_), .B(_11158__bF_buf4), .C(_11196_), .Y(_11197_) );
	OAI21X1 OAI21X1_4426 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(_11127__bF_buf4), .C(biu_pc_9_), .Y(_11198_) );
	OAI21X1 OAI21X1_4427 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11197_), .C(_11198_), .Y(csr_gpr_iu_csr_tval_9_) );
	INVX1 INVX1_1791 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_10_), .Y(_11199_) );
	OAI21X1 OAI21X1_4428 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11199_), .C(_11158__bF_buf3), .Y(_11200_) );
	OAI21X1 OAI21X1_4429 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_11158__bF_buf2), .C(_11200_), .Y(_11201_) );
	OAI21X1 OAI21X1_4430 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11127__bF_buf3), .C(biu_pc_10_), .Y(_11202_) );
	OAI21X1 OAI21X1_4431 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11201_), .C(_11202_), .Y(csr_gpr_iu_csr_tval_10_) );
	INVX1 INVX1_1792 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_11_), .Y(_11203_) );
	OAI21X1 OAI21X1_4432 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11203_), .C(_11158__bF_buf1), .Y(_11204_) );
	OAI21X1 OAI21X1_4433 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_11_), .B(_11158__bF_buf0), .C(_11204_), .Y(_11205_) );
	OAI21X1 OAI21X1_4434 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(_11127__bF_buf2), .C(biu_pc_11_), .Y(_11206_) );
	OAI21X1 OAI21X1_4435 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11205_), .C(_11206_), .Y(csr_gpr_iu_csr_tval_11_) );
	INVX1 INVX1_1793 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_12_), .Y(_11207_) );
	OAI21X1 OAI21X1_4436 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11207_), .C(_11158__bF_buf7), .Y(_11208_) );
	OAI21X1 OAI21X1_4437 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_11158__bF_buf6), .C(_11208_), .Y(_11209_) );
	OAI21X1 OAI21X1_4438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf1), .C(biu_pc_12_), .Y(_11210_) );
	OAI21X1 OAI21X1_4439 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11209_), .C(_11210_), .Y(csr_gpr_iu_csr_tval_12_) );
	INVX1 INVX1_1794 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_13_), .Y(_11211_) );
	OAI21X1 OAI21X1_4440 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11211_), .C(_11158__bF_buf5), .Y(_11212_) );
	OAI21X1 OAI21X1_4441 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_13_bF_buf3), .B(_11158__bF_buf4), .C(_11212_), .Y(_11213_) );
	OAI21X1 OAI21X1_4442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf0), .C(biu_pc_13_), .Y(_11214_) );
	OAI21X1 OAI21X1_4443 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11213_), .C(_11214_), .Y(csr_gpr_iu_csr_tval_13_) );
	INVX1 INVX1_1795 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_14_), .Y(_11215_) );
	OAI21X1 OAI21X1_4444 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11215_), .C(_11158__bF_buf3), .Y(_11216_) );
	OAI21X1 OAI21X1_4445 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_11158__bF_buf2), .C(_11216_), .Y(_11217_) );
	OAI21X1 OAI21X1_4446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(_11127__bF_buf4), .C(biu_pc_14_), .Y(_11218_) );
	OAI21X1 OAI21X1_4447 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11217_), .C(_11218_), .Y(csr_gpr_iu_csr_tval_14_) );
	INVX1 INVX1_1796 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf5), .Y(_11219_) );
	OAI21X1 OAI21X1_4448 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11219_), .C(_11158__bF_buf1), .Y(_11220_) );
	OAI21X1 OAI21X1_4449 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_15_bF_buf0), .B(_11158__bF_buf0), .C(_11220_), .Y(_11221_) );
	OAI21X1 OAI21X1_4450 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(_11127__bF_buf3), .C(biu_pc_15_), .Y(_11222_) );
	OAI21X1 OAI21X1_4451 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11221_), .C(_11222_), .Y(csr_gpr_iu_csr_tval_15_) );
	INVX1 INVX1_1797 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_16_), .Y(_11223_) );
	OAI21X1 OAI21X1_4452 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11223_), .C(_11158__bF_buf7), .Y(_11224_) );
	OAI21X1 OAI21X1_4453 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_11158__bF_buf6), .C(_11224_), .Y(_11225_) );
	OAI21X1 OAI21X1_4454 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11127__bF_buf2), .C(biu_pc_16_), .Y(_11226_) );
	OAI21X1 OAI21X1_4455 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11225_), .C(_11226_), .Y(csr_gpr_iu_csr_tval_16_) );
	INVX1 INVX1_1798 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_17_), .Y(_11227_) );
	OAI21X1 OAI21X1_4456 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11227_), .C(_11158__bF_buf5), .Y(_11228_) );
	OAI21X1 OAI21X1_4457 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_17_bF_buf0), .B(_11158__bF_buf4), .C(_11228_), .Y(_11229_) );
	OAI21X1 OAI21X1_4458 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(_11127__bF_buf1), .C(biu_pc_17_), .Y(_11230_) );
	OAI21X1 OAI21X1_4459 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11229_), .C(_11230_), .Y(csr_gpr_iu_csr_tval_17_) );
	INVX1 INVX1_1799 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .Y(_11231_) );
	OAI21X1 OAI21X1_4460 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11231_), .C(_11158__bF_buf3), .Y(_11232_) );
	OAI21X1 OAI21X1_4461 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_11158__bF_buf2), .C(_11232_), .Y(_11233_) );
	OAI21X1 OAI21X1_4462 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf0), .C(biu_pc_18_), .Y(_11234_) );
	OAI21X1 OAI21X1_4463 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11233_), .C(_11234_), .Y(csr_gpr_iu_csr_tval_18_) );
	INVX1 INVX1_1800 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_19_), .Y(_11235_) );
	OAI21X1 OAI21X1_4464 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11235_), .C(_11158__bF_buf1), .Y(_11236_) );
	OAI21X1 OAI21X1_4465 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_19_bF_buf1), .B(_11158__bF_buf0), .C(_11236_), .Y(_11237_) );
	OAI21X1 OAI21X1_4466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf4), .C(biu_pc_19_), .Y(_11238_) );
	OAI21X1 OAI21X1_4467 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11237_), .C(_11238_), .Y(csr_gpr_iu_csr_tval_19_) );
	INVX1 INVX1_1801 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf5), .Y(_11239_) );
	OAI21X1 OAI21X1_4468 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11239_), .C(_11158__bF_buf7), .Y(_11240_) );
	OAI21X1 OAI21X1_4469 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_11158__bF_buf6), .C(_11240_), .Y(_11241_) );
	OAI21X1 OAI21X1_4470 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(_11127__bF_buf3), .C(biu_pc_20_), .Y(_11242_) );
	OAI21X1 OAI21X1_4471 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11241_), .C(_11242_), .Y(csr_gpr_iu_csr_tval_20_) );
	INVX1 INVX1_1802 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf1), .Y(_11243_) );
	OAI21X1 OAI21X1_4472 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11243_), .C(_11158__bF_buf5), .Y(_11244_) );
	OAI21X1 OAI21X1_4473 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_21_bF_buf2), .B(_11158__bF_buf4), .C(_11244_), .Y(_11245_) );
	OAI21X1 OAI21X1_4474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(_11127__bF_buf2), .C(biu_pc_21_), .Y(_11246_) );
	OAI21X1 OAI21X1_4475 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11245_), .C(_11246_), .Y(csr_gpr_iu_csr_tval_21_) );
	INVX1 INVX1_1803 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf3), .Y(_11247_) );
	OAI21X1 OAI21X1_4476 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11247_), .C(_11158__bF_buf3), .Y(_11248_) );
	OAI21X1 OAI21X1_4477 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_11158__bF_buf2), .C(_11248_), .Y(_11249_) );
	OAI21X1 OAI21X1_4478 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11127__bF_buf1), .C(biu_pc_22_), .Y(_11250_) );
	OAI21X1 OAI21X1_4479 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11249_), .C(_11250_), .Y(csr_gpr_iu_csr_tval_22_) );
	INVX1 INVX1_1804 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .Y(_11251_) );
	OAI21X1 OAI21X1_4480 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11251_), .C(_11158__bF_buf1), .Y(_11252_) );
	OAI21X1 OAI21X1_4481 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_23_bF_buf0), .B(_11158__bF_buf0), .C(_11252_), .Y(_11253_) );
	OAI21X1 OAI21X1_4482 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(_11127__bF_buf0), .C(biu_pc_23_), .Y(_11254_) );
	OAI21X1 OAI21X1_4483 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11253_), .C(_11254_), .Y(csr_gpr_iu_csr_tval_23_) );
	INVX1 INVX1_1805 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_11255_) );
	OAI21X1 OAI21X1_4484 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11255_), .C(_11158__bF_buf7), .Y(_11256_) );
	OAI21X1 OAI21X1_4485 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_11158__bF_buf6), .C(_11256_), .Y(_11257_) );
	OAI21X1 OAI21X1_4486 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf4), .C(biu_pc_24_), .Y(_11258_) );
	OAI21X1 OAI21X1_4487 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11257_), .C(_11258_), .Y(csr_gpr_iu_csr_tval_24_) );
	INVX1 INVX1_1806 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf2), .Y(_11259_) );
	OAI21X1 OAI21X1_4488 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11259_), .C(_11158__bF_buf5), .Y(_11260_) );
	OAI21X1 OAI21X1_4489 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_25_bF_buf2), .B(_11158__bF_buf4), .C(_11260_), .Y(_11261_) );
	OAI21X1 OAI21X1_4490 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf3), .C(biu_pc_25_), .Y(_11262_) );
	OAI21X1 OAI21X1_4491 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11261_), .C(_11262_), .Y(csr_gpr_iu_csr_tval_25_) );
	INVX1 INVX1_1807 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf0), .Y(_11263_) );
	OAI21X1 OAI21X1_4492 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11263_), .C(_11158__bF_buf3), .Y(_11264_) );
	OAI21X1 OAI21X1_4493 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .B(_11158__bF_buf2), .C(_11264_), .Y(_11265_) );
	OAI21X1 OAI21X1_4494 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf4), .B(_11127__bF_buf2), .C(biu_pc_26_), .Y(_11266_) );
	OAI21X1 OAI21X1_4495 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11265_), .C(_11266_), .Y(csr_gpr_iu_csr_tval_26_) );
	INVX1 INVX1_1808 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf2), .Y(_11267_) );
	OAI21X1 OAI21X1_4496 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf1), .B(_11267_), .C(_11158__bF_buf1), .Y(_11268_) );
	OAI21X1 OAI21X1_4497 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_27_bF_buf3), .B(_11158__bF_buf0), .C(_11268_), .Y(_11269_) );
	OAI21X1 OAI21X1_4498 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf3), .B(_11127__bF_buf1), .C(biu_pc_27_), .Y(_11270_) );
	OAI21X1 OAI21X1_4499 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf2), .B(_11269_), .C(_11270_), .Y(csr_gpr_iu_csr_tval_27_) );
	INVX1 INVX1_1809 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf3), .Y(_11271_) );
	OAI21X1 OAI21X1_4500 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf0), .B(_11271_), .C(_11158__bF_buf7), .Y(_11272_) );
	OAI21X1 OAI21X1_4501 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_11158__bF_buf6), .C(_11272_), .Y(_11273_) );
	OAI21X1 OAI21X1_4502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf2), .B(_11127__bF_buf0), .C(biu_pc_28_), .Y(_11274_) );
	OAI21X1 OAI21X1_4503 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf1), .B(_11273_), .C(_11274_), .Y(csr_gpr_iu_csr_tval_28_) );
	INVX1 INVX1_1810 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf0), .Y(_11275_) );
	OAI21X1 OAI21X1_4504 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf4), .B(_11275_), .C(_11158__bF_buf5), .Y(_11276_) );
	OAI21X1 OAI21X1_4505 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_29_bF_buf2), .B(_11158__bF_buf4), .C(_11276_), .Y(_11277_) );
	OAI21X1 OAI21X1_4506 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf1), .B(_11127__bF_buf4), .C(biu_pc_29_), .Y(_11278_) );
	OAI21X1 OAI21X1_4507 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf0), .B(_11277_), .C(_11278_), .Y(csr_gpr_iu_csr_tval_29_) );
	INVX1 INVX1_1811 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf1), .Y(_11279_) );
	OAI21X1 OAI21X1_4508 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf3), .B(_11279_), .C(_11158__bF_buf3), .Y(_11280_) );
	OAI21X1 OAI21X1_4509 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_11158__bF_buf2), .C(_11280_), .Y(_11281_) );
	OAI21X1 OAI21X1_4510 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf0), .B(_11127__bF_buf3), .C(biu_pc_30_), .Y(_11282_) );
	OAI21X1 OAI21X1_4511 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf4), .B(_11281_), .C(_11282_), .Y(csr_gpr_iu_csr_tval_30_) );
	INVX1 INVX1_1812 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .Y(_11283_) );
	OAI21X1 OAI21X1_4512 ( .gnd(gnd), .vdd(vdd), .A(_11119__bF_buf2), .B(_11283_), .C(_11158__bF_buf1), .Y(_11284_) );
	OAI21X1 OAI21X1_4513 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_31_bF_buf0), .B(_11158__bF_buf0), .C(_11284_), .Y(_11285_) );
	OAI21X1 OAI21X1_4514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_page_fault_bF_buf5), .B(_11127__bF_buf2), .C(biu_pc_31_), .Y(_11286_) );
	OAI21X1 OAI21X1_4515 ( .gnd(gnd), .vdd(vdd), .A(_11156__bF_buf3), .B(_11285_), .C(_11286_), .Y(csr_gpr_iu_csr_tval_31_) );
	NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_10988_), .B(_10987_), .Y(_11287_) );
	INVX1 INVX1_1813 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf17), .Y(_11288_) );
	OAI21X1 OAI21X1_4516 ( .gnd(gnd), .vdd(vdd), .A(ext_int), .B(_11287_), .C(_11288_), .Y(_11289_) );
	AOI21X1 AOI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_11016_), .B(_11287_), .C(_11289_), .Y(_10983_) );
	OAI21X1 OAI21X1_4517 ( .gnd(gnd), .vdd(vdd), .A(soft_int), .B(_11287_), .C(_11288_), .Y(_11290_) );
	AOI21X1 AOI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_11024_), .B(_11287_), .C(_11290_), .Y(_10984_) );
	OAI21X1 OAI21X1_4518 ( .gnd(gnd), .vdd(vdd), .A(timer_int), .B(_11287_), .C(_11288_), .Y(_11291_) );
	AOI21X1 AOI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .B(_11287_), .C(_11291_), .Y(_10985_) );
	DFFPOSX1 DFFPOSX1_1908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_10985_), .Q(csr_gpr_iu_int_ctrl_timer_int) );
	DFFPOSX1 DFFPOSX1_1909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_10984_), .Q(csr_gpr_iu_int_ctrl_soft_int) );
	DFFPOSX1 DFFPOSX1_1910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_10983_), .Q(csr_gpr_iu_int_ctrl_ext_int) );
	NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_0_), .B(exu_alu_shift_counter_1_), .Y(_13387_) );
	INVX1 INVX1_1814 ( .gnd(gnd), .vdd(vdd), .A(_13387_), .Y(_13388_) );
	NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_2_), .B(_13388_), .Y(_13389_) );
	NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_3_), .B(exu_alu_shift_counter_4_), .Y(_13390_) );
	NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_13390_), .B(_13389_), .Y(_13391_) );
	INVX8 INVX8_93 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf7), .Y(_13392_) );
	INVX1 INVX1_1815 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .Y(_13393_) );
	NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_1_), .B(_13393_), .Y(_13394_) );
	INVX1 INVX1_1816 ( .gnd(gnd), .vdd(vdd), .A(_13394_), .Y(_13395_) );
	NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(_13395_), .Y(_13396_) );
	INVX8 INVX8_94 ( .gnd(gnd), .vdd(vdd), .A(_13396_), .Y(_13397_) );
	NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .B(_13397__bF_buf4), .Y(_13398_) );
	INVX1 INVX1_1817 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_slli), .Y(_13399_) );
	NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_srli), .B(csr_gpr_iu_ins_dec_srai), .Y(_13400_) );
	NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_13399_), .B(_13400_), .Y(_13401_) );
	INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .Y(_13402_) );
	INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .Y(_13403_) );
	INVX1 INVX1_1818 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sllp), .Y(_13404_) );
	NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_srlp), .B(csr_gpr_iu_ins_dec_srap), .Y(_13405_) );
	NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_13404_), .B(_13405_), .Y(_13406_) );
	INVX1 INVX1_1819 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .Y(_13407_) );
	OAI21X1 OAI21X1_4519 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13407_), .C(_13402_), .Y(_13408_) );
	OAI21X1 OAI21X1_4520 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf4), .B(_13402_), .C(_13408_), .Y(_13409_) );
	NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_13409_), .B(_13398__bF_buf6), .Y(_13410_) );
	OAI21X1 OAI21X1_4521 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_0_), .B(_13398__bF_buf5), .C(_13410_), .Y(_13411_) );
	INVX8 INVX8_95 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf16), .Y(_13412_) );
	INVX1 INVX1_1820 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_0_), .Y(_13413_) );
	NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_slli), .B(csr_gpr_iu_ins_dec_sllp), .Y(_13414_) );
	INVX8 INVX8_96 ( .gnd(gnd), .vdd(vdd), .A(_13414_), .Y(_13415_) );
	NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_13400_), .B(_13405_), .Y(_13416_) );
	NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf6), .B(_13416__bF_buf4), .Y(_13417_) );
	INVX1 INVX1_1821 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .Y(_13418_) );
	NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_13413_), .B(_13418_), .Y(_13419_) );
	OAI21X1 OAI21X1_4522 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_0_), .B(_13417_), .C(_13391__bF_buf6), .Y(_13420_) );
	OAI21X1 OAI21X1_4523 ( .gnd(gnd), .vdd(vdd), .A(_13420_), .B(_13419_), .C(_13412__bF_buf4), .Y(_13421_) );
	AOI21X1 AOI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_13411_), .B(_13392__bF_buf7), .C(_13421_), .Y(_11294__0_) );
	NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_13388_), .B(_13417_), .Y(_13422_) );
	INVX1 INVX1_1822 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_1_), .Y(_13423_) );
	AOI21X1 AOI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_13418_), .B(_13413_), .C(_13423_), .Y(_13424_) );
	OAI21X1 OAI21X1_4524 ( .gnd(gnd), .vdd(vdd), .A(_13422_), .B(_13424_), .C(_13391__bF_buf5), .Y(_13425_) );
	NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(_13407_), .Y(_13426_) );
	AOI22X1 AOI22X1_647 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_21_bF_buf0), .B(_13401_), .C(csr_gpr_iu_rs2_1_), .D(_13426_), .Y(_13427_) );
	AOI21X1 AOI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf4), .B(_13427_), .C(_13391__bF_buf4), .Y(_13428_) );
	OAI21X1 OAI21X1_4525 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_1_), .B(_13398__bF_buf3), .C(_13428_), .Y(_13429_) );
	AOI21X1 AOI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_13429_), .B(_13425_), .C(rst_bF_buf15), .Y(_11294__1_) );
	OAI21X1 OAI21X1_4526 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf5), .B(_13416__bF_buf3), .C(_13389_), .Y(_13430_) );
	INVX1 INVX1_1823 ( .gnd(gnd), .vdd(vdd), .A(_13430_), .Y(_13431_) );
	INVX1 INVX1_1824 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_2_), .Y(_13432_) );
	NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_13432_), .B(_13422_), .Y(_13433_) );
	OAI21X1 OAI21X1_4527 ( .gnd(gnd), .vdd(vdd), .A(_13431_), .B(_13433_), .C(_13391__bF_buf3), .Y(_13434_) );
	INVX4 INVX4_33 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .Y(_13435_) );
	INVX1 INVX1_1825 ( .gnd(gnd), .vdd(vdd), .A(_13426_), .Y(_13436_) );
	NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf2), .B(_13401_), .Y(_13437_) );
	OAI21X1 OAI21X1_4528 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13436_), .C(_13437_), .Y(_13438_) );
	INVX1 INVX1_1826 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .Y(_13439_) );
	NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf2), .B(_13397__bF_buf3), .Y(_13440_) );
	NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .B(_13440_), .Y(_13441_) );
	INVX1 INVX1_1827 ( .gnd(gnd), .vdd(vdd), .A(_13441__bF_buf4), .Y(_13442_) );
	NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_13438_), .B(_13442_), .Y(_13443_) );
	AOI21X1 AOI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13434_), .C(rst_bF_buf14), .Y(_11294__2_) );
	XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_13430_), .B(exu_alu_shift_counter_3_), .Y(_13444_) );
	NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .B(_13398__bF_buf2), .Y(_13445_) );
	NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_23_), .B(_13401_), .C(_13398__bF_buf1), .Y(_13446_) );
	OAI21X1 OAI21X1_4529 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .B(_13445_), .C(_13446_), .Y(_13447_) );
	OAI21X1 OAI21X1_4530 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf1), .B(_13447_), .C(_13412__bF_buf3), .Y(_13448_) );
	AOI21X1 AOI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf0), .B(_13444_), .C(_13448_), .Y(_11294__3_) );
	OAI21X1 OAI21X1_4531 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_3_), .B(_13430_), .C(exu_alu_shift_counter_4_), .Y(_13449_) );
	INVX1 INVX1_1828 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_13450_) );
	INVX4 INVX4_34 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_4_), .Y(_13451_) );
	OAI22X1 OAI22X1_817 ( .gnd(gnd), .vdd(vdd), .A(_13450_), .B(_13402_), .C(_13451_), .D(_13436_), .Y(_13452_) );
	NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_13452_), .B(_13442_), .Y(_13453_) );
	AOI21X1 AOI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_13453_), .B(_13449_), .C(rst_bF_buf13), .Y(_11294__4_) );
	NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .B(_13397__bF_buf2), .Y(_13454_) );
	INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .Y(_13455_) );
	NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(amominu), .B(amomin), .Y(_13456_) );
	NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(amomaxu), .B(amomax), .Y(_13457_) );
	NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .B(_13457_), .Y(_13458_) );
	INVX8 INVX8_97 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf8), .Y(_13459_) );
	NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(amoswap), .Y(_13460_) );
	NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(amoxor_bF_buf3), .C(amoor), .Y(_13461_) );
	AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_13461_), .B(_13460_), .Y(_13462_) );
	NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf4), .B(_13462__bF_buf3), .Y(_13463_) );
	INVX8 INVX8_98 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf2), .Y(_13464_) );
	NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(amoor), .Y(_13465_) );
	NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_13464__bF_buf3), .B(_13460_), .C(_13465_), .Y(_13466_) );
	OAI21X1 OAI21X1_4532 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf6), .C(biu_biu_data_out_0_), .Y(_13467_) );
	OAI21X1 OAI21X1_4533 ( .gnd(gnd), .vdd(vdd), .A(_13455_), .B(_13463__bF_buf4), .C(_13467_), .Y(_13468_) );
	INVX1 INVX1_1829 ( .gnd(gnd), .vdd(vdd), .A(_13468_), .Y(_13469_) );
	NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf1), .B(csr_gpr_iu_ins_dec_xorp), .Y(_13470_) );
	INVX4 INVX4_35 ( .gnd(gnd), .vdd(vdd), .A(_13470__bF_buf4), .Y(_13471_) );
	OAI21X1 OAI21X1_4534 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf0), .B(csr_gpr_iu_ins_dec_xorp), .C(_13403_), .Y(_13472_) );
	OAI21X1 OAI21X1_4535 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(_13471_), .C(_13472_), .Y(_13473_) );
	AOI21X1 AOI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .B(_13473_), .C(_13464__bF_buf2), .Y(_13474_) );
	OAI21X1 OAI21X1_4536 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .B(_13473_), .C(_13474_), .Y(_13475_) );
	NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf5), .Y(_13476_) );
	NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .B(_13476__bF_buf3), .Y(_13477_) );
	NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(addp_bF_buf4), .Y(_13478_) );
	INVX1 INVX1_1830 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .Y(_13479_) );
	NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(addi_bF_buf6), .Y(_13480_) );
	OAI21X1 OAI21X1_4537 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(_13479_), .C(_13480_), .Y(_13481_) );
	NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_13478__bF_buf4), .B(_13481_), .Y(_13482_) );
	OAI21X1 OAI21X1_4538 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(addp_bF_buf3), .C(csr_gpr_iu_rs2_0_), .Y(_13483_) );
	AOI22X1 AOI22X1_648 ( .gnd(gnd), .vdd(vdd), .A(_13482_), .B(_13483_), .C(_13467_), .D(_13477_), .Y(_13484_) );
	OAI21X1 OAI21X1_4539 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13478__bF_buf3), .C(_13482_), .Y(_13485_) );
	NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_13485_), .B(_13468_), .Y(_13486_) );
	NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .B(_13486_), .Y(_13487_) );
	NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf0), .B(amoand), .Y(_13488_) );
	INVX4 INVX4_36 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf3), .Y(_13489_) );
	AOI22X1 AOI22X1_649 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(amoswap), .C(_13489_), .D(_13487_), .Y(_13490_) );
	NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(_13490_), .Y(_13491_) );
	INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_0_), .Y(_13492_) );
	INVX1 INVX1_1831 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_28_), .Y(_13493_) );
	INVX4 INVX4_37 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .Y(_13494_) );
	NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_29_), .B(_13494_), .Y(_13495_) );
	OAI21X1 OAI21X1_4540 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_13493_), .C(_13495_), .Y(_13496_) );
	INVX4 INVX4_38 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .Y(_13497_) );
	NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_30_), .B(_13497_), .Y(_13498_) );
	INVX1 INVX1_1832 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_30_), .Y(_13499_) );
	XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(biu_biu_data_out_31_), .Y(_13500_) );
	OAI21X1 OAI21X1_4541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_13499_), .C(_13500_), .Y(_13501_) );
	NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(_13501_), .Y(_13502_) );
	NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_13493_), .Y(_13503_) );
	OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(biu_biu_data_out_29_), .Y(_13504_) );
	NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_13503_), .B(_13504_), .C(_13502_), .Y(_13505_) );
	OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .B(_13496_), .Y(_13506_) );
	INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_26_), .Y(_13507_) );
	INVX4 INVX4_39 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_27_), .Y(_13508_) );
	NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_27_), .B(_13508_), .Y(_13509_) );
	INVX1 INVX1_1833 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_27_), .Y(_13510_) );
	NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_27_), .B(_13510_), .Y(_13511_) );
	NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_13509_), .B(_13511_), .Y(_13512_) );
	OAI21X1 OAI21X1_4542 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_13507_), .C(_13512_), .Y(_13513_) );
	AOI21X1 AOI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_13507_), .C(_13513_), .Y(_13514_) );
	INVX4 INVX4_40 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .Y(_13515_) );
	INVX4 INVX4_41 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .Y(_13516_) );
	NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_24_), .B(_13516_), .Y(_13517_) );
	AOI21X1 AOI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(biu_biu_data_out_25_), .C(_13517_), .Y(_13518_) );
	INVX1 INVX1_1834 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_25_), .Y(_13519_) );
	AOI22X1 AOI22X1_650 ( .gnd(gnd), .vdd(vdd), .A(_13519_), .B(csr_gpr_iu_rs2_25_), .C(_13516_), .D(biu_biu_data_out_24_), .Y(_13520_) );
	NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_13518_), .B(_13520_), .C(_13514_), .Y(_13521_) );
	OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .B(_13521_), .Y(_13522_) );
	INVX1 INVX1_1835 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_21_), .Y(_13523_) );
	INVX1 INVX1_1836 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_20_), .Y(_13524_) );
	OAI22X1 OAI22X1_818 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_13523_), .C(csr_gpr_iu_rs2_20_), .D(_13524_), .Y(_13525_) );
	INVX4 INVX4_42 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_23_), .Y(_13526_) );
	NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_23_), .B(_13526_), .Y(_13527_) );
	INVX1 INVX1_1837 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_23_), .Y(_13528_) );
	NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_23_), .B(_13528_), .Y(_13529_) );
	OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .B(_13529_), .Y(_13530_) );
	INVX1 INVX1_1838 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_22_), .Y(_13531_) );
	NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_13531_), .Y(_13532_) );
	INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .Y(_13533_) );
	NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_22_), .B(_13533_), .Y(_13534_) );
	NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_13532_), .B(_13534_), .Y(_13535_) );
	NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_13535_), .B(_13530_), .Y(_13536_) );
	INVX1 INVX1_1839 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .Y(_13537_) );
	INVX4 INVX4_43 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .Y(_13538_) );
	NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_13523_), .Y(_13539_) );
	OAI21X1 OAI21X1_4543 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(biu_biu_data_out_20_), .C(_13539_), .Y(_13540_) );
	OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .B(_13540_), .Y(_13541_) );
	NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_13525_), .B(_13541_), .Y(_13542_) );
	INVX1 INVX1_1840 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_18_), .Y(_13543_) );
	NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_13543_), .Y(_13544_) );
	INVX4 INVX4_44 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .Y(_13545_) );
	NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_19_), .B(_13545_), .Y(_13546_) );
	INVX1 INVX1_1841 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_19_), .Y(_13547_) );
	NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_13547_), .Y(_13548_) );
	NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_13546_), .B(_13548_), .Y(_13549_) );
	INVX4 INVX4_45 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .Y(_13550_) );
	NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_18_), .B(_13550_), .Y(_13551_) );
	NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .B(_13551_), .C(_13549_), .Y(_13552_) );
	INVX1 INVX1_1842 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_17_), .Y(_13553_) );
	INVX1 INVX1_1843 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_16_), .Y(_13554_) );
	AOI22X1 AOI22X1_651 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .B(csr_gpr_iu_rs2_17_), .C(csr_gpr_iu_rs2_16_), .D(_13554_), .Y(_13555_) );
	INVX4 INVX4_46 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .Y(_13556_) );
	NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_13553_), .Y(_13557_) );
	AOI21X1 AOI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(biu_biu_data_out_16_), .C(_13557_), .Y(_13558_) );
	NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_13555_), .B(_13558_), .Y(_13559_) );
	NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_13559_), .B(_13552_), .Y(_13560_) );
	NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_13560_), .B(_13542_), .Y(_13561_) );
	NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_13522_), .B(_13561_), .Y(_13562_) );
	INVX1 INVX1_1844 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_13_), .Y(_13563_) );
	INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .Y(_13564_) );
	NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_12_), .B(_13564_), .Y(_13565_) );
	OAI21X1 OAI21X1_4544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_13563_), .C(_13565_), .Y(_13566_) );
	INVX1 INVX1_1845 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_14_), .Y(_13567_) );
	NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_13567_), .Y(_13568_) );
	INVX1 INVX1_1846 ( .gnd(gnd), .vdd(vdd), .A(_13568_), .Y(_13569_) );
	INVX4 INVX4_47 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .Y(_13570_) );
	NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .B(_13570_), .Y(_13571_) );
	INVX1 INVX1_1847 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .Y(_13572_) );
	NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_13572_), .Y(_13573_) );
	NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_13571_), .B(_13573_), .Y(_13574_) );
	OAI21X1 OAI21X1_4545 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_13567_), .C(_13574_), .Y(_13575_) );
	NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .B(_13575_), .Y(_13576_) );
	INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .Y(_13577_) );
	NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_13_), .B(_13577_), .Y(_13578_) );
	INVX1 INVX1_1848 ( .gnd(gnd), .vdd(vdd), .A(_13578_), .Y(_13579_) );
	INVX1 INVX1_1849 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_12_), .Y(_13580_) );
	NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_13580_), .Y(_13581_) );
	NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(_13579_), .B(_13581_), .C(_13576_), .Y(_13582_) );
	NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_13566_), .B(_13582_), .Y(_13583_) );
	INVX1 INVX1_1850 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_10_), .Y(_13584_) );
	NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_10_), .B(_13584_), .Y(_13585_) );
	INVX1 INVX1_1851 ( .gnd(gnd), .vdd(vdd), .A(_13585_), .Y(_13586_) );
	INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .Y(_13587_) );
	NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_11_), .B(_13587_), .Y(_13588_) );
	INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_11_), .Y(_13589_) );
	NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_13589_), .Y(_13590_) );
	NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_13588_), .B(_13590_), .Y(_13591_) );
	OAI21X1 OAI21X1_4546 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_10_), .B(_13584_), .C(_13591_), .Y(_13592_) );
	OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_13592_), .B(_13586_), .Y(_13593_) );
	INVX1 INVX1_1852 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_9_), .Y(_13594_) );
	NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .B(_13594_), .Y(_13595_) );
	INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .Y(_13596_) );
	NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_9_), .B(_13596_), .Y(_13597_) );
	NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_13595_), .B(_13597_), .Y(_13598_) );
	INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_8_), .Y(_13599_) );
	NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .B(_13599_), .Y(_13600_) );
	NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .B(_13599_), .Y(_13601_) );
	INVX1 INVX1_1853 ( .gnd(gnd), .vdd(vdd), .A(_13601_), .Y(_13602_) );
	NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_13600_), .B(_13602_), .C(_13598_), .Y(_13603_) );
	NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_13603_), .B(_13593_), .Y(_13604_) );
	NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13583_), .Y(_13605_) );
	INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_6_), .Y(_13606_) );
	NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .B(_13606_), .Y(_13607_) );
	INVX1 INVX1_1854 ( .gnd(gnd), .vdd(vdd), .A(_13607_), .Y(_13608_) );
	XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(biu_biu_data_out_7_bF_buf0), .Y(_13609_) );
	OAI21X1 OAI21X1_4547 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .B(_13606_), .C(_13609_), .Y(_13610_) );
	OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_13610_), .B(_13608_), .Y(_13611_) );
	INVX4 INVX4_48 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_5_), .Y(_13612_) );
	NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_5_), .B(_13612_), .Y(_13613_) );
	NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .B(_13451_), .Y(_13614_) );
	NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .B(_13451_), .Y(_13615_) );
	NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_5_), .B(_13612_), .Y(_13616_) );
	NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .B(_13616_), .Y(_13617_) );
	NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(_13613_), .B(_13614_), .C(_13617_), .Y(_13618_) );
	NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .B(_13611_), .Y(_13619_) );
	NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_2_), .B(_13435_), .Y(_13620_) );
	INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_2_), .Y(_13621_) );
	INVX4 INVX4_49 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .Y(_13622_) );
	NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .B(_13622_), .Y(_13623_) );
	INVX1 INVX1_1855 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .Y(_13624_) );
	NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .B(_13624_), .Y(_13625_) );
	NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_13623_), .B(_13625_), .Y(_13626_) );
	OAI21X1 OAI21X1_4548 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .B(_13621_), .C(_13626_), .Y(_13627_) );
	OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_13627_), .B(_13620_), .Y(_13628_) );
	INVX1 INVX1_1856 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_1_), .Y(_13629_) );
	INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .Y(_13630_) );
	NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(_13629_), .Y(_13631_) );
	OAI21X1 OAI21X1_4549 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_13492_), .C(_13631_), .Y(_13632_) );
	AOI21X1 AOI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(biu_biu_data_out_1_), .C(_13632_), .Y(_13633_) );
	AOI21X1 AOI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(_13629_), .C(_13633_), .Y(_13634_) );
	AOI21X1 AOI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13620_), .C(_13623_), .Y(_13635_) );
	OAI21X1 OAI21X1_4550 ( .gnd(gnd), .vdd(vdd), .A(_13634_), .B(_13628_), .C(_13635_), .Y(_13636_) );
	NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_13636_), .Y(_13637_) );
	AOI21X1 AOI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .B(_13613_), .C(_13616_), .Y(_13638_) );
	NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_13638_), .B(_13611_), .Y(_13639_) );
	INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .Y(_13640_) );
	INVX1 INVX1_1857 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_7_bF_buf3), .Y(_13641_) );
	OAI21X1 OAI21X1_4551 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(_13641_), .C(_13608_), .Y(_13642_) );
	OAI21X1 OAI21X1_4552 ( .gnd(gnd), .vdd(vdd), .A(_13640_), .B(biu_biu_data_out_7_bF_buf2), .C(_13642_), .Y(_13643_) );
	NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_13643_), .B(_13639_), .Y(_13644_) );
	AOI21X1 AOI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_13637_), .B(_13644_), .C(_13605_), .Y(_13645_) );
	AOI21X1 AOI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_13598_), .B(_13601_), .C(_13597_), .Y(_13646_) );
	AOI21X1 AOI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_13591_), .B(_13586_), .C(_13588_), .Y(_13647_) );
	OAI21X1 OAI21X1_4553 ( .gnd(gnd), .vdd(vdd), .A(_13646_), .B(_13593_), .C(_13647_), .Y(_13648_) );
	NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_13648_), .B(_13583_), .Y(_13649_) );
	AOI21X1 AOI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(biu_biu_data_out_13_), .C(_13581_), .Y(_13650_) );
	OAI21X1 OAI21X1_4554 ( .gnd(gnd), .vdd(vdd), .A(_13578_), .B(_13650_), .C(_13576_), .Y(_13651_) );
	AOI21X1 AOI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_13574_), .B(_13569_), .C(_13571_), .Y(_13652_) );
	NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(_13651_), .B(_13652_), .C(_13649_), .Y(_13653_) );
	OAI21X1 OAI21X1_4555 ( .gnd(gnd), .vdd(vdd), .A(_13653_), .B(_13645_), .C(_13562_), .Y(_13654_) );
	INVX1 INVX1_1858 ( .gnd(gnd), .vdd(vdd), .A(_13546_), .Y(_13655_) );
	OAI21X1 OAI21X1_4556 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .B(_13548_), .C(_13655_), .Y(_13656_) );
	OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_13555_), .B(_13557_), .Y(_13657_) );
	NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13552_), .Y(_13658_) );
	OAI21X1 OAI21X1_4557 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .B(_13658_), .C(_13542_), .Y(_13659_) );
	INVX1 INVX1_1859 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .Y(_13660_) );
	OAI21X1 OAI21X1_4558 ( .gnd(gnd), .vdd(vdd), .A(_13532_), .B(_13529_), .C(_13660_), .Y(_13661_) );
	NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_13523_), .Y(_13662_) );
	NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(_13524_), .Y(_13663_) );
	OAI21X1 OAI21X1_4559 ( .gnd(gnd), .vdd(vdd), .A(_13663_), .B(_13662_), .C(_13539_), .Y(_13664_) );
	AOI21X1 AOI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .B(_13664_), .C(_13661_), .Y(_13665_) );
	AOI21X1 AOI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_13659_), .B(_13665_), .C(_13522_), .Y(_13666_) );
	OAI21X1 OAI21X1_4560 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_13519_), .C(_13517_), .Y(_13667_) );
	OAI21X1 OAI21X1_4561 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(biu_biu_data_out_25_), .C(_13667_), .Y(_13668_) );
	NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_13507_), .C(_13512_), .Y(_13669_) );
	OAI21X1 OAI21X1_4562 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(biu_biu_data_out_27_), .C(_13669_), .Y(_13670_) );
	AOI21X1 AOI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_13514_), .B(_13668_), .C(_13670_), .Y(_13671_) );
	INVX1 INVX1_1860 ( .gnd(gnd), .vdd(vdd), .A(_13495_), .Y(_13672_) );
	OAI21X1 OAI21X1_4563 ( .gnd(gnd), .vdd(vdd), .A(_13503_), .B(_13672_), .C(_13504_), .Y(_13673_) );
	INVX4 INVX4_50 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .Y(_13674_) );
	INVX1 INVX1_1861 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_31_), .Y(_13675_) );
	OAI21X1 OAI21X1_4564 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_13675_), .C(_13498_), .Y(_13676_) );
	OAI21X1 OAI21X1_4565 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(biu_biu_data_out_31_), .C(_13676_), .Y(_13677_) );
	AOI21X1 AOI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(_13673_), .C(_13677_), .Y(_13678_) );
	OAI21X1 OAI21X1_4566 ( .gnd(gnd), .vdd(vdd), .A(_13671_), .B(_13506_), .C(_13678_), .Y(_13679_) );
	NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_13679_), .B(_13666_), .Y(_13680_) );
	NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_13654_), .B(_13680_), .Y(_13681_) );
	AOI21X1 AOI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_13492_), .C(_13628_), .Y(_13682_) );
	NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_13633_), .B(_13682_), .C(_13619_), .Y(_13683_) );
	NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_13683_), .B(_13605_), .Y(_13684_) );
	AOI21X1 AOI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_13562_), .B(_13684_), .C(_13457_), .Y(_13685_) );
	NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .B(_13681_), .Y(_13686_) );
	AOI21X1 AOI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .B(_13685_), .C(_13686_), .Y(_13687_) );
	OAI21X1 OAI21X1_4567 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_13687__bF_buf7), .C(_13458__bF_buf5), .Y(_13688_) );
	AOI21X1 AOI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_13492_), .B(_13687__bF_buf6), .C(_13688_), .Y(_13689_) );
	OAI21X1 OAI21X1_4568 ( .gnd(gnd), .vdd(vdd), .A(_13491_), .B(_13689_), .C(_13454__bF_buf4), .Y(_13690_) );
	INVX1 INVX1_1862 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sc_w), .Y(_13691_) );
	INVX1 INVX1_1863 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_2_), .Y(_13692_) );
	OAI21X1 OAI21X1_4569 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_0_), .B(biu_exce_chk_opc_1_), .C(_13692_), .Y(_13693_) );
	NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_13691_), .B(_13693_), .Y(_13694_) );
	INVX8 INVX8_99 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf0), .Y(_13695_) );
	NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13695__bF_buf5), .Y(_13696_) );
	INVX1 INVX1_1864 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_0_), .Y(_13697_) );
	OAI21X1 OAI21X1_4570 ( .gnd(gnd), .vdd(vdd), .A(_13697_), .B(_13396_), .C(_13392__bF_buf6), .Y(_13698_) );
	AOI21X1 AOI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_13696_), .B(_13694__bF_buf4), .C(_13698_), .Y(_13699_) );
	OAI21X1 OAI21X1_4571 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_0_), .B(_13392__bF_buf5), .C(_13412__bF_buf2), .Y(_13700_) );
	AOI21X1 AOI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_13690_), .B(_13699_), .C(_13700_), .Y(_11293__0_) );
	NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_13629_), .B(_13687__bF_buf5), .Y(_13701_) );
	OAI21X1 OAI21X1_4572 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(_13687__bF_buf4), .C(_13701_), .Y(_13702_) );
	NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf3), .B(_13702_), .Y(_13703_) );
	OAI21X1 OAI21X1_4573 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf4), .C(_13629_), .Y(_13704_) );
	INVX1 INVX1_1865 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_1_), .Y(_13705_) );
	NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_13705_), .B(_13459__bF_buf2), .C(_13462__bF_buf2), .Y(_13706_) );
	OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(addp_bF_buf2), .Y(_13707_) );
	INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_1_), .Y(_13708_) );
	NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(_13708_), .Y(_13709_) );
	OAI21X1 OAI21X1_4574 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(biu_pc_1_), .C(_13709_), .Y(_13710_) );
	OAI21X1 OAI21X1_4575 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(addp_bF_buf1), .C(csr_gpr_iu_rs2_1_), .Y(_13711_) );
	OAI21X1 OAI21X1_4576 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13710_), .C(_13711_), .Y(_13712_) );
	NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .B(_13712_), .C(_13706_), .Y(_13713_) );
	OAI21X1 OAI21X1_4577 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf3), .C(biu_biu_data_out_1_), .Y(_13714_) );
	NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_1_), .B(_13476__bF_buf2), .Y(_13715_) );
	INVX1 INVX1_1866 ( .gnd(gnd), .vdd(vdd), .A(_13712_), .Y(_13716_) );
	NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(_13714_), .B(_13715_), .C(_13716_), .Y(_13717_) );
	NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_13713_), .B(_13717_), .Y(_13718_) );
	XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_13718_), .B(_13484_), .Y(_13719_) );
	OAI21X1 OAI21X1_4578 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(amoand), .C(_13719_), .Y(_13720_) );
	OAI21X1 OAI21X1_4579 ( .gnd(gnd), .vdd(vdd), .A(_13705_), .B(_13463__bF_buf3), .C(_13714_), .Y(_13721_) );
	OAI21X1 OAI21X1_4580 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf3), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_1_), .Y(_13722_) );
	OAI21X1 OAI21X1_4581 ( .gnd(gnd), .vdd(vdd), .A(_13708_), .B(_13471_), .C(_13722_), .Y(_13723_) );
	AOI21X1 AOI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .B(_13723_), .C(_13464__bF_buf1), .Y(_13724_) );
	OAI21X1 OAI21X1_4582 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .B(_13723_), .C(_13724_), .Y(_13725_) );
	INVX4 INVX4_51 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf3), .Y(_13726_) );
	AOI21X1 AOI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(amoswap), .C(_13726_), .Y(_13727_) );
	NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(_13725_), .B(_13727_), .C(_13720_), .Y(_13728_) );
	INVX1 INVX1_1867 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_1_), .Y(_13729_) );
	AOI21X1 AOI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_13729_), .B(_13397__bF_buf1), .C(_13398__bF_buf6), .Y(_13730_) );
	OAI21X1 OAI21X1_4583 ( .gnd(gnd), .vdd(vdd), .A(_13728_), .B(_13703_), .C(_13730_), .Y(_13731_) );
	NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(_13695__bF_buf4), .Y(_13732_) );
	AOI21X1 AOI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_13732_), .B(_13694__bF_buf3), .C(_13391__bF_buf7), .Y(_13733_) );
	OAI21X1 OAI21X1_4584 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_1_), .B(_13392__bF_buf4), .C(_13412__bF_buf1), .Y(_13734_) );
	AOI21X1 AOI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_13731_), .B(_13733_), .C(_13734_), .Y(_11293__1_) );
	NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .B(_13459__bF_buf1), .C(_13462__bF_buf1), .Y(_13735_) );
	OAI21X1 OAI21X1_4585 ( .gnd(gnd), .vdd(vdd), .A(_13621_), .B(_13476__bF_buf1), .C(_13735_), .Y(_13736_) );
	NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .B(_13470__bF_buf3), .Y(_13737_) );
	OAI21X1 OAI21X1_4586 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13470__bF_buf2), .C(_13737_), .Y(_13738_) );
	OAI21X1 OAI21X1_4587 ( .gnd(gnd), .vdd(vdd), .A(_13738_), .B(_13736_), .C(amoxor_bF_buf2), .Y(_13739_) );
	AOI21X1 AOI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_13736_), .B(_13738_), .C(_13739_), .Y(_13740_) );
	AOI21X1 AOI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .B(amoswap), .C(_13740_), .Y(_13741_) );
	OAI21X1 OAI21X1_4588 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf2), .B(_13466__bF_buf2), .C(_13492_), .Y(_13742_) );
	NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_13455_), .B(_13459__bF_buf0), .C(_13462__bF_buf0), .Y(_13743_) );
	NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(_13742_), .B(_13485_), .C(_13743_), .Y(_13744_) );
	OAI21X1 OAI21X1_4589 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf0), .B(addp_bF_buf0), .C(_13630_), .Y(_13745_) );
	NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_13478__bF_buf2), .B(_13710_), .Y(_13746_) );
	AOI22X1 AOI22X1_652 ( .gnd(gnd), .vdd(vdd), .A(_13745_), .B(_13746_), .C(_13704_), .D(_13706_), .Y(_13747_) );
	OAI21X1 OAI21X1_4590 ( .gnd(gnd), .vdd(vdd), .A(_13744_), .B(_13747_), .C(_13713_), .Y(_13748_) );
	OAI21X1 OAI21X1_4591 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf1), .C(biu_biu_data_out_2_), .Y(_13749_) );
	INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .Y(_13750_) );
	NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(csr_gpr_iu_imm12_2_), .Y(_13751_) );
	OAI21X1 OAI21X1_4592 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(_13750_), .C(_13751_), .Y(_13752_) );
	OAI21X1 OAI21X1_4593 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(addp_bF_buf4), .C(_13435_), .Y(_13753_) );
	OAI21X1 OAI21X1_4594 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13752_), .C(_13753_), .Y(_13754_) );
	INVX1 INVX1_1868 ( .gnd(gnd), .vdd(vdd), .A(_13754_), .Y(_13755_) );
	NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13755_), .C(_13735_), .Y(_13756_) );
	OAI21X1 OAI21X1_4595 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf0), .C(_13621_), .Y(_13757_) );
	INVX1 INVX1_1869 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .Y(_13758_) );
	NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_13758_), .B(_13459__bF_buf4), .C(_13462__bF_buf3), .Y(_13759_) );
	NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_13757_), .B(_13754_), .C(_13759_), .Y(_13760_) );
	NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_13760_), .B(_13756_), .Y(_13761_) );
	XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_13748_), .B(_13761_), .Y(_13762_) );
	INVX1 INVX1_1870 ( .gnd(gnd), .vdd(vdd), .A(_13762_), .Y(_13763_) );
	OAI21X1 OAI21X1_4596 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf2), .B(_13763_), .C(_13741_), .Y(_13764_) );
	OAI21X1 OAI21X1_4597 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .B(_13687__bF_buf3), .C(_13458__bF_buf8), .Y(_13765_) );
	AOI21X1 AOI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_13621_), .B(_13687__bF_buf2), .C(_13765_), .Y(_13766_) );
	OAI21X1 OAI21X1_4598 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_13766_), .C(_13454__bF_buf2), .Y(_13767_) );
	NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13695__bF_buf3), .Y(_13768_) );
	INVX1 INVX1_1871 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_2_), .Y(_13769_) );
	OAI21X1 OAI21X1_4599 ( .gnd(gnd), .vdd(vdd), .A(_13769_), .B(_13396_), .C(_13392__bF_buf3), .Y(_13770_) );
	AOI21X1 AOI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_13768_), .B(_13694__bF_buf2), .C(_13770_), .Y(_13771_) );
	OAI21X1 OAI21X1_4600 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_2_), .B(_13392__bF_buf2), .C(_13412__bF_buf0), .Y(_13772_) );
	AOI21X1 AOI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_13767_), .B(_13771_), .C(_13772_), .Y(_11293__2_) );
	OAI21X1 OAI21X1_4601 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf6), .B(_13397__bF_buf0), .C(biu_biu_data_in_3_), .Y(_13773_) );
	INVX1 INVX1_1872 ( .gnd(gnd), .vdd(vdd), .A(_13694__bF_buf1), .Y(_13774_) );
	NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_13774_), .B(_13445_), .Y(_13775_) );
	INVX8 INVX8_100 ( .gnd(gnd), .vdd(vdd), .A(amoswap), .Y(_13776_) );
	INVX1 INVX1_1873 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .Y(_13777_) );
	NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_13459__bF_buf3), .C(_13462__bF_buf2), .Y(_13778_) );
	OAI21X1 OAI21X1_4602 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .B(_13476__bF_buf0), .C(_13778_), .Y(_13779_) );
	OAI21X1 OAI21X1_4603 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf1), .B(csr_gpr_iu_ins_dec_xorp), .C(_13622_), .Y(_13780_) );
	OAI21X1 OAI21X1_4604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_3_), .B(_13471_), .C(_13780_), .Y(_13781_) );
	AOI21X1 AOI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_13779_), .B(_13781_), .C(_13464__bF_buf0), .Y(_13782_) );
	OAI21X1 OAI21X1_4605 ( .gnd(gnd), .vdd(vdd), .A(_13779_), .B(_13781_), .C(_13782_), .Y(_13783_) );
	OAI21X1 OAI21X1_4606 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_13776__bF_buf3), .C(_13783_), .Y(_13784_) );
	OAI21X1 OAI21X1_4607 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf6), .C(biu_biu_data_out_3_), .Y(_13785_) );
	NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .B(_13459__bF_buf2), .C(_13462__bF_buf1), .Y(_13786_) );
	INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .Y(_13787_) );
	NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(csr_gpr_iu_imm12_3_), .Y(_13788_) );
	OAI21X1 OAI21X1_4608 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(_13787_), .C(_13788_), .Y(_13789_) );
	OAI21X1 OAI21X1_4609 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(addp_bF_buf3), .C(_13622_), .Y(_13790_) );
	OAI21X1 OAI21X1_4610 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13789_), .C(_13790_), .Y(_13791_) );
	INVX1 INVX1_1874 ( .gnd(gnd), .vdd(vdd), .A(_13791_), .Y(_13792_) );
	NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_13785_), .B(_13792_), .C(_13786_), .Y(_13793_) );
	OAI21X1 OAI21X1_4611 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf5), .C(_13624_), .Y(_13794_) );
	NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_13794_), .B(_13791_), .C(_13778_), .Y(_13795_) );
	NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_13795_), .B(_13793_), .Y(_13796_) );
	NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(_13757_), .B(_13755_), .C(_13759_), .Y(_13797_) );
	INVX1 INVX1_1875 ( .gnd(gnd), .vdd(vdd), .A(_13797_), .Y(_13798_) );
	AOI21X1 AOI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_13748_), .B(_13761_), .C(_13798_), .Y(_13799_) );
	XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_13799_), .B(_13796_), .Y(_13800_) );
	AOI21X1 AOI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_13800_), .B(_13489_), .C(_13784_), .Y(_13801_) );
	NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_3_), .B(_13687__bF_buf1), .Y(_13802_) );
	OAI21X1 OAI21X1_4612 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_13687__bF_buf0), .C(_13802_), .Y(_13803_) );
	NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf5), .B(_13803_), .Y(_13804_) );
	AOI21X1 AOI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_13804_), .B(_13801_), .C(_13726_), .Y(_13805_) );
	OAI21X1 OAI21X1_4613 ( .gnd(gnd), .vdd(vdd), .A(_13775_), .B(_13805_), .C(_13392__bF_buf1), .Y(_13806_) );
	AOI21X1 AOI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_13806_), .B(_13773_), .C(rst_bF_buf12), .Y(_11293__3_) );
	OAI21X1 OAI21X1_4614 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf5), .B(_13397__bF_buf4), .C(biu_biu_data_in_4_), .Y(_13807_) );
	NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_4_), .B(_13398__bF_buf5), .Y(_13808_) );
	NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_13774_), .B(_13808_), .Y(_13809_) );
	INVX1 INVX1_1876 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_4_), .Y(_13810_) );
	NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_13810_), .B(_13459__bF_buf1), .C(_13462__bF_buf0), .Y(_13811_) );
	OAI21X1 OAI21X1_4615 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .B(_13476__bF_buf3), .C(_13811_), .Y(_13812_) );
	INVX1 INVX1_1877 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_4_), .Y(_13813_) );
	OAI21X1 OAI21X1_4616 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf0), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_4_), .Y(_13814_) );
	OAI21X1 OAI21X1_4617 ( .gnd(gnd), .vdd(vdd), .A(_13813_), .B(_13471_), .C(_13814_), .Y(_13815_) );
	AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_13812_), .B(_13815_), .Y(_13816_) );
	NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_13815_), .B(_13812_), .Y(_13817_) );
	OAI21X1 OAI21X1_4618 ( .gnd(gnd), .vdd(vdd), .A(_13817_), .B(_13816_), .C(amoxor_bF_buf3), .Y(_13818_) );
	NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .B(_13687__bF_buf7), .Y(_13819_) );
	OAI21X1 OAI21X1_4619 ( .gnd(gnd), .vdd(vdd), .A(_13451_), .B(_13687__bF_buf6), .C(_13819_), .Y(_13820_) );
	AOI22X1 AOI22X1_653 ( .gnd(gnd), .vdd(vdd), .A(_13756_), .B(_13760_), .C(_13793_), .D(_13795_), .Y(_13821_) );
	NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(_13794_), .B(_13792_), .C(_13778_), .Y(_13822_) );
	AOI21X1 AOI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_13778_), .B(_13794_), .C(_13792_), .Y(_13823_) );
	OAI21X1 OAI21X1_4620 ( .gnd(gnd), .vdd(vdd), .A(_13797_), .B(_13823_), .C(_13822_), .Y(_13824_) );
	AOI21X1 AOI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_13821_), .B(_13748_), .C(_13824_), .Y(_13825_) );
	OAI21X1 OAI21X1_4621 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf4), .C(biu_biu_data_out_4_), .Y(_13826_) );
	NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_4_), .B(_13459__bF_buf0), .C(_13462__bF_buf3), .Y(_13827_) );
	INVX1 INVX1_1878 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_4_), .Y(_13828_) );
	NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(csr_gpr_iu_imm12_4_), .Y(_13829_) );
	OAI21X1 OAI21X1_4622 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(_13828_), .C(_13829_), .Y(_13830_) );
	OAI21X1 OAI21X1_4623 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(addp_bF_buf2), .C(_13451_), .Y(_13831_) );
	OAI21X1 OAI21X1_4624 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13830_), .C(_13831_), .Y(_13832_) );
	INVX1 INVX1_1879 ( .gnd(gnd), .vdd(vdd), .A(_13832_), .Y(_13833_) );
	NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(_13826_), .B(_13833_), .C(_13827_), .Y(_13834_) );
	INVX1 INVX1_1880 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_4_), .Y(_13835_) );
	OAI21X1 OAI21X1_4625 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf3), .C(_13835_), .Y(_13836_) );
	NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_13836_), .B(_13832_), .C(_13811_), .Y(_13837_) );
	NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_13837_), .B(_13834_), .Y(_13838_) );
	INVX1 INVX1_1881 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .Y(_13839_) );
	NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_13839_), .B(_13825_), .Y(_13840_) );
	NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_13748_), .B(_13821_), .Y(_13841_) );
	INVX1 INVX1_1882 ( .gnd(gnd), .vdd(vdd), .A(_13824_), .Y(_13842_) );
	NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_13842_), .B(_13841_), .Y(_13843_) );
	NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .B(_13843_), .Y(_13844_) );
	NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_13844_), .Y(_13845_) );
	OAI21X1 OAI21X1_4626 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf0), .B(amoand), .C(_13845_), .Y(_13846_) );
	OAI21X1 OAI21X1_4627 ( .gnd(gnd), .vdd(vdd), .A(_13451_), .B(_13776__bF_buf2), .C(_13846_), .Y(_13847_) );
	AOI21X1 AOI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_13820_), .B(_13458__bF_buf2), .C(_13847_), .Y(_13848_) );
	AOI21X1 AOI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_13848_), .B(_13818_), .C(_13726_), .Y(_13849_) );
	OAI21X1 OAI21X1_4628 ( .gnd(gnd), .vdd(vdd), .A(_13809_), .B(_13849_), .C(_13392__bF_buf0), .Y(_13850_) );
	AOI21X1 AOI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_13850_), .B(_13807_), .C(rst_bF_buf11), .Y(_11293__4_) );
	INVX1 INVX1_1883 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_5_), .Y(_13851_) );
	NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_13851_), .B(_13687__bF_buf5), .Y(_13852_) );
	OAI21X1 OAI21X1_4629 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_5_), .B(_13687__bF_buf4), .C(_13852_), .Y(_13853_) );
	INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .Y(_13854_) );
	OAI21X1 OAI21X1_4630 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf2), .C(biu_biu_data_out_5_), .Y(_13855_) );
	OAI21X1 OAI21X1_4631 ( .gnd(gnd), .vdd(vdd), .A(_13854_), .B(_13463__bF_buf2), .C(_13855_), .Y(_13856_) );
	NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf1), .B(_13470__bF_buf1), .Y(_13857_) );
	OAI21X1 OAI21X1_4632 ( .gnd(gnd), .vdd(vdd), .A(_13612_), .B(_13470__bF_buf0), .C(_13857_), .Y(_13858_) );
	OAI21X1 OAI21X1_4633 ( .gnd(gnd), .vdd(vdd), .A(_13858_), .B(_13856_), .C(amoxor_bF_buf2), .Y(_13859_) );
	AOI21X1 AOI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_13856_), .B(_13858_), .C(_13859_), .Y(_13860_) );
	AOI21X1 AOI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_5_), .B(amoswap), .C(_13860_), .Y(_13861_) );
	OAI21X1 OAI21X1_4634 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf4), .B(_13853_), .C(_13861_), .Y(_13862_) );
	INVX1 INVX1_1884 ( .gnd(gnd), .vdd(vdd), .A(_13812_), .Y(_13863_) );
	AOI21X1 AOI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_13863_), .B(_13833_), .C(_13840_), .Y(_13864_) );
	OAI21X1 OAI21X1_4635 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf1), .C(_13851_), .Y(_13865_) );
	NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_13854_), .B(_13476__bF_buf2), .Y(_13866_) );
	INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .Y(_13867_) );
	NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(biu_ins_25_bF_buf0), .Y(_13868_) );
	OAI21X1 OAI21X1_4636 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(_13867_), .C(_13868_), .Y(_13869_) );
	OAI21X1 OAI21X1_4637 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(addp_bF_buf1), .C(_13612_), .Y(_13870_) );
	OAI21X1 OAI21X1_4638 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13869_), .C(_13870_), .Y(_13871_) );
	INVX1 INVX1_1885 ( .gnd(gnd), .vdd(vdd), .A(_13871_), .Y(_13872_) );
	NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(_13865_), .B(_13872_), .C(_13866_), .Y(_13873_) );
	NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .B(_13476__bF_buf1), .Y(_13874_) );
	NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_13871_), .C(_13874_), .Y(_13875_) );
	NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_13873_), .B(_13875_), .Y(_13876_) );
	XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_13864_), .B(_13876_), .Y(_13877_) );
	OAI21X1 OAI21X1_4639 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf1), .B(_13877_), .C(_13454__bF_buf1), .Y(_13878_) );
	INVX1 INVX1_1886 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_5_), .Y(_13879_) );
	AOI21X1 AOI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_13879_), .B(_13397__bF_buf3), .C(_13398__bF_buf4), .Y(_13880_) );
	OAI21X1 OAI21X1_4640 ( .gnd(gnd), .vdd(vdd), .A(_13878_), .B(_13862_), .C(_13880_), .Y(_13881_) );
	NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_13612_), .B(_13695__bF_buf2), .Y(_13882_) );
	AOI21X1 AOI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_13882_), .B(_13694__bF_buf0), .C(_13391__bF_buf4), .Y(_13883_) );
	OAI21X1 OAI21X1_4641 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_5_), .B(_13392__bF_buf7), .C(_13412__bF_buf4), .Y(_13884_) );
	AOI21X1 AOI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_13883_), .C(_13884_), .Y(_11293__5_) );
	INVX4 INVX4_52 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .Y(_13885_) );
	NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_6_), .B(_13687__bF_buf3), .Y(_13886_) );
	OAI21X1 OAI21X1_4642 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_13687__bF_buf2), .C(_13886_), .Y(_13887_) );
	NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf8), .B(_13887_), .Y(_13888_) );
	NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .B(_13459__bF_buf3), .C(_13462__bF_buf2), .Y(_13889_) );
	OAI21X1 OAI21X1_4643 ( .gnd(gnd), .vdd(vdd), .A(_13606_), .B(_13476__bF_buf0), .C(_13889_), .Y(_13890_) );
	NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf3), .B(_13470__bF_buf4), .Y(_13891_) );
	OAI21X1 OAI21X1_4644 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_13470__bF_buf3), .C(_13891_), .Y(_13892_) );
	OAI21X1 OAI21X1_4645 ( .gnd(gnd), .vdd(vdd), .A(_13892_), .B(_13890_), .C(amoxor_bF_buf1), .Y(_13893_) );
	AOI21X1 AOI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_13890_), .B(_13892_), .C(_13893_), .Y(_13894_) );
	AOI21X1 AOI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .B(amoswap), .C(_13894_), .Y(_13895_) );
	OAI21X1 OAI21X1_4646 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf0), .C(biu_biu_data_out_6_), .Y(_13896_) );
	INVX1 INVX1_1887 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_6_), .Y(_13897_) );
	NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(biu_ins_26_bF_buf2), .Y(_13898_) );
	OAI21X1 OAI21X1_4647 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(_13897_), .C(_13898_), .Y(_13899_) );
	OAI21X1 OAI21X1_4648 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(addp_bF_buf0), .C(_13885_), .Y(_13900_) );
	OAI21X1 OAI21X1_4649 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13899_), .C(_13900_), .Y(_13901_) );
	INVX1 INVX1_1888 ( .gnd(gnd), .vdd(vdd), .A(_13901_), .Y(_13902_) );
	NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(_13896_), .B(_13902_), .C(_13889_), .Y(_13903_) );
	OAI21X1 OAI21X1_4650 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf6), .C(_13606_), .Y(_13904_) );
	INVX1 INVX1_1889 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .Y(_13905_) );
	NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(_13905_), .B(_13459__bF_buf2), .C(_13462__bF_buf1), .Y(_13906_) );
	NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(_13904_), .B(_13901_), .C(_13906_), .Y(_13907_) );
	NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_13907_), .B(_13903_), .Y(_13908_) );
	OAI21X1 OAI21X1_4651 ( .gnd(gnd), .vdd(vdd), .A(_13812_), .B(_13832_), .C(_13873_), .Y(_13909_) );
	OAI21X1 OAI21X1_4652 ( .gnd(gnd), .vdd(vdd), .A(_13909_), .B(_13840_), .C(_13875_), .Y(_13910_) );
	XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_13910_), .B(_13908_), .Y(_13911_) );
	AOI21X1 AOI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_13911_), .B(_13489_), .C(_13726_), .Y(_13912_) );
	NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(_13895_), .B(_13912_), .C(_13888_), .Y(_13913_) );
	INVX1 INVX1_1890 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_6_), .Y(_13914_) );
	AOI21X1 AOI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_13914_), .B(_13397__bF_buf2), .C(_13398__bF_buf3), .Y(_13915_) );
	NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_13915_), .B(_13913_), .Y(_13916_) );
	NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_13695__bF_buf1), .Y(_13917_) );
	AOI21X1 AOI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_13917_), .B(_13694__bF_buf4), .C(_13391__bF_buf3), .Y(_13918_) );
	OAI21X1 OAI21X1_4653 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_6_), .B(_13392__bF_buf6), .C(_13412__bF_buf3), .Y(_13919_) );
	AOI21X1 AOI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_13916_), .B(_13918_), .C(_13919_), .Y(_11293__6_) );
	OAI21X1 OAI21X1_4654 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_6_), .B(_13476__bF_buf3), .C(_13906_), .Y(_13920_) );
	NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_13901_), .B(_13920_), .Y(_13921_) );
	INVX1 INVX1_1891 ( .gnd(gnd), .vdd(vdd), .A(_13921_), .Y(_13922_) );
	INVX1 INVX1_1892 ( .gnd(gnd), .vdd(vdd), .A(_13908_), .Y(_13923_) );
	OAI21X1 OAI21X1_4655 ( .gnd(gnd), .vdd(vdd), .A(_13923_), .B(_13910_), .C(_13922_), .Y(_13924_) );
	OAI21X1 OAI21X1_4656 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf5), .B(_13466__bF_buf5), .C(biu_biu_data_out_7_bF_buf1), .Y(_13925_) );
	INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(_13925_), .Y(_13926_) );
	INVX1 INVX1_1893 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_7_), .Y(_13927_) );
	NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_13927_), .B(_13458__bF_buf4), .C(_13466__bF_buf4), .Y(_13928_) );
	INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .Y(_13929_) );
	NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(biu_ins_27_bF_buf1), .Y(_13930_) );
	OAI21X1 OAI21X1_4657 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(_13929_), .C(_13930_), .Y(_13931_) );
	OAI21X1 OAI21X1_4658 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(addp_bF_buf4), .C(_13640_), .Y(_13932_) );
	OAI21X1 OAI21X1_4659 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13931_), .C(_13932_), .Y(_13933_) );
	INVX1 INVX1_1894 ( .gnd(gnd), .vdd(vdd), .A(_13933_), .Y(_13934_) );
	OAI21X1 OAI21X1_4660 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .B(_13926_), .C(_13934_), .Y(_13935_) );
	INVX1 INVX1_1895 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .Y(_13936_) );
	NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_13925_), .B(_13933_), .C(_13936_), .Y(_13937_) );
	NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_13935_), .B(_13937_), .Y(_13938_) );
	XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_13924_), .B(_13938_), .Y(_13939_) );
	NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf0), .B(_13939_), .Y(_13940_) );
	NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_13641_), .B(_13687__bF_buf1), .Y(_13941_) );
	OAI21X1 OAI21X1_4661 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(_13687__bF_buf0), .C(_13941_), .Y(_13942_) );
	NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .B(_13926_), .Y(_13943_) );
	INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(_13943_), .Y(_13944_) );
	INVX1 INVX1_1896 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf0), .Y(_13945_) );
	OAI21X1 OAI21X1_4662 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf0), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_7_), .Y(_13946_) );
	OAI21X1 OAI21X1_4663 ( .gnd(gnd), .vdd(vdd), .A(_13945_), .B(_13471_), .C(_13946_), .Y(_13947_) );
	OAI21X1 OAI21X1_4664 ( .gnd(gnd), .vdd(vdd), .A(_13947_), .B(_13944_), .C(amoxor_bF_buf3), .Y(_13948_) );
	AOI21X1 AOI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_13947_), .C(_13948_), .Y(_13949_) );
	OAI21X1 OAI21X1_4665 ( .gnd(gnd), .vdd(vdd), .A(_13640_), .B(_13776__bF_buf1), .C(_13454__bF_buf0), .Y(_13950_) );
	NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_13950_), .B(_13949_), .Y(_13951_) );
	OAI21X1 OAI21X1_4666 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf1), .B(_13942_), .C(_13951_), .Y(_13952_) );
	INVX1 INVX1_1897 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_7_), .Y(_13953_) );
	AOI21X1 AOI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_13953_), .B(_13397__bF_buf1), .C(_13398__bF_buf2), .Y(_13954_) );
	OAI21X1 OAI21X1_4667 ( .gnd(gnd), .vdd(vdd), .A(_13940_), .B(_13952_), .C(_13954_), .Y(_13955_) );
	NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_13640_), .B(_13695__bF_buf0), .Y(_13956_) );
	AOI21X1 AOI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_13956_), .B(_13694__bF_buf3), .C(_13391__bF_buf2), .Y(_13957_) );
	OAI21X1 OAI21X1_4668 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_7_), .B(_13392__bF_buf5), .C(_13412__bF_buf2), .Y(_13958_) );
	AOI21X1 AOI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_13955_), .B(_13957_), .C(_13958_), .Y(_11293__7_) );
	NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .B(_13687__bF_buf7), .Y(_13959_) );
	OAI21X1 OAI21X1_4669 ( .gnd(gnd), .vdd(vdd), .A(_13599_), .B(_13687__bF_buf6), .C(_13959_), .Y(_13960_) );
	NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13960_), .Y(_13961_) );
	INVX1 INVX1_1898 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_8_), .Y(_13962_) );
	NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .B(_13459__bF_buf0), .C(_13462__bF_buf0), .Y(_13963_) );
	OAI21X1 OAI21X1_4670 ( .gnd(gnd), .vdd(vdd), .A(_13962_), .B(_13476__bF_buf2), .C(_13963_), .Y(_13964_) );
	INVX1 INVX1_1899 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf2), .Y(_13965_) );
	OAI21X1 OAI21X1_4671 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf2), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_8_), .Y(_13966_) );
	OAI21X1 OAI21X1_4672 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13471_), .C(_13966_), .Y(_13967_) );
	OAI21X1 OAI21X1_4673 ( .gnd(gnd), .vdd(vdd), .A(_13967_), .B(_13964_), .C(amoxor_bF_buf1), .Y(_13968_) );
	AOI21X1 AOI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(_13967_), .C(_13968_), .Y(_13969_) );
	AOI21X1 AOI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_8_), .B(amoswap), .C(_13969_), .Y(_13970_) );
	NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(_13873_), .B(_13875_), .C(_13838_), .Y(_13971_) );
	NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(_13935_), .B(_13937_), .C(_13908_), .Y(_13972_) );
	NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_13971_), .B(_13972_), .Y(_13973_) );
	OAI21X1 OAI21X1_4674 ( .gnd(gnd), .vdd(vdd), .A(_13856_), .B(_13872_), .C(_13909_), .Y(_13974_) );
	OAI21X1 OAI21X1_4675 ( .gnd(gnd), .vdd(vdd), .A(_13920_), .B(_13901_), .C(_13935_), .Y(_13975_) );
	OAI21X1 OAI21X1_4676 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_13934_), .C(_13975_), .Y(_13976_) );
	OAI21X1 OAI21X1_4677 ( .gnd(gnd), .vdd(vdd), .A(_13972_), .B(_13974_), .C(_13976_), .Y(_13977_) );
	AOI21X1 AOI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_13843_), .B(_13973_), .C(_13977_), .Y(_13978_) );
	OAI21X1 OAI21X1_4678 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf2), .B(_13466__bF_buf3), .C(_13962_), .Y(_13979_) );
	INVX1 INVX1_1900 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .Y(_13980_) );
	NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13459__bF_buf4), .C(_13462__bF_buf3), .Y(_13981_) );
	INVX1 INVX1_1901 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_8_), .Y(_13982_) );
	NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(biu_ins_28_bF_buf1), .Y(_13983_) );
	OAI21X1 OAI21X1_4679 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(_13982_), .C(_13983_), .Y(_13984_) );
	OAI21X1 OAI21X1_4680 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf0), .B(addp_bF_buf3), .C(_13599_), .Y(_11295_) );
	OAI21X1 OAI21X1_4681 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13984_), .C(_11295_), .Y(_11296_) );
	INVX1 INVX1_1902 ( .gnd(gnd), .vdd(vdd), .A(_11296_), .Y(_11297_) );
	NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(_13979_), .B(_11297_), .C(_13981_), .Y(_11298_) );
	OAI21X1 OAI21X1_4682 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf2), .C(biu_biu_data_out_8_), .Y(_11299_) );
	NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_11299_), .B(_11296_), .C(_13963_), .Y(_11300_) );
	AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_11298_), .B(_11300_), .Y(_11301_) );
	XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_13978_), .B(_11301_), .Y(_11302_) );
	AOI21X1 AOI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_11302_), .B(_13489_), .C(_13726_), .Y(_11303_) );
	NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(_13970_), .B(_11303_), .C(_13961_), .Y(_11304_) );
	INVX1 INVX1_1903 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_8_), .Y(_11305_) );
	AOI21X1 AOI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_11305_), .B(_13397__bF_buf0), .C(_13398__bF_buf1), .Y(_11306_) );
	NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_11306_), .B(_11304_), .Y(_11307_) );
	NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_13599_), .B(_13695__bF_buf5), .Y(_11308_) );
	AOI21X1 AOI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_13694__bF_buf2), .C(_13391__bF_buf1), .Y(_11309_) );
	OAI21X1 OAI21X1_4683 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_8_), .B(_13392__bF_buf4), .C(_13412__bF_buf1), .Y(_11310_) );
	AOI21X1 AOI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_11307_), .B(_11309_), .C(_11310_), .Y(_11293__8_) );
	NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_11300_), .B(_11298_), .Y(_11311_) );
	OAI21X1 OAI21X1_4684 ( .gnd(gnd), .vdd(vdd), .A(_11311_), .B(_13978_), .C(_11298_), .Y(_11312_) );
	OAI21X1 OAI21X1_4685 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf1), .C(biu_biu_data_out_9_), .Y(_11313_) );
	NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_9_), .B(_13476__bF_buf1), .Y(_11314_) );
	INVX1 INVX1_1904 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .Y(_11315_) );
	NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(biu_ins_29_bF_buf3), .Y(_11316_) );
	OAI21X1 OAI21X1_4686 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(_11315_), .C(_11316_), .Y(_11317_) );
	OAI21X1 OAI21X1_4687 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(addp_bF_buf2), .C(_13596_), .Y(_11318_) );
	OAI21X1 OAI21X1_4688 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_11317_), .C(_11318_), .Y(_11319_) );
	AOI21X1 AOI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_11314_), .B(_11313_), .C(_11319_), .Y(_11320_) );
	INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(_11313_), .Y(_11321_) );
	INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_9_), .Y(_11322_) );
	NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_11322_), .B(_13458__bF_buf8), .C(_13466__bF_buf0), .Y(_11323_) );
	INVX1 INVX1_1905 ( .gnd(gnd), .vdd(vdd), .A(_11319_), .Y(_11324_) );
	NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .B(_11324_), .C(_11321_), .Y(_11325_) );
	NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11325_), .Y(_11326_) );
	XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_11312_), .B(_11326_), .Y(_11327_) );
	OAI21X1 OAI21X1_4689 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(amoand), .C(_11327_), .Y(_11328_) );
	NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_9_), .B(_13687__bF_buf5), .Y(_11329_) );
	OAI21X1 OAI21X1_4690 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .B(_13687__bF_buf4), .C(_11329_), .Y(_11330_) );
	NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_11330_), .Y(_11331_) );
	OAI21X1 OAI21X1_4691 ( .gnd(gnd), .vdd(vdd), .A(_11322_), .B(_13463__bF_buf1), .C(_11313_), .Y(_11332_) );
	INVX1 INVX1_1906 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf2), .Y(_11333_) );
	OAI21X1 OAI21X1_4692 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf0), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_9_), .Y(_11334_) );
	OAI21X1 OAI21X1_4693 ( .gnd(gnd), .vdd(vdd), .A(_11333_), .B(_13471_), .C(_11334_), .Y(_11335_) );
	OAI21X1 OAI21X1_4694 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11332_), .C(amoxor_bF_buf3), .Y(_11336_) );
	AOI21X1 AOI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_11332_), .B(_11335_), .C(_11336_), .Y(_11337_) );
	AOI21X1 AOI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .B(amoswap), .C(_11337_), .Y(_11338_) );
	NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(_11328_), .B(_11338_), .C(_11331_), .Y(_11339_) );
	INVX1 INVX1_1907 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_9_), .Y(_11340_) );
	AOI21X1 AOI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_11340_), .B(_13397__bF_buf4), .C(_13398__bF_buf0), .Y(_11341_) );
	OAI21X1 OAI21X1_4695 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_11339_), .C(_11341_), .Y(_11342_) );
	NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .B(_13695__bF_buf4), .Y(_11343_) );
	AOI21X1 AOI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_11343_), .B(_13694__bF_buf1), .C(_13391__bF_buf0), .Y(_11344_) );
	OAI21X1 OAI21X1_4696 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_9_), .B(_13392__bF_buf3), .C(_13412__bF_buf0), .Y(_11345_) );
	AOI21X1 AOI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_11342_), .B(_11344_), .C(_11345_), .Y(_11293__9_) );
	OAI21X1 OAI21X1_4697 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf6), .C(biu_biu_data_out_10_), .Y(_11346_) );
	NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .B(_13476__bF_buf0), .Y(_11347_) );
	INVX1 INVX1_1908 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf0), .Y(_11348_) );
	NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(biu_pc_10_), .Y(_11349_) );
	AOI21X1 AOI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(_11348_), .C(_11349_), .Y(_11350_) );
	INVX4 INVX4_53 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_10_), .Y(_11351_) );
	OAI21X1 OAI21X1_4698 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(addp_bF_buf1), .C(_11351_), .Y(_11352_) );
	OAI21X1 OAI21X1_4699 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_11350_), .C(_11352_), .Y(_11353_) );
	AOI21X1 AOI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_11347_), .B(_11346_), .C(_11353_), .Y(_11354_) );
	AOI21X1 AOI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_13462__bF_buf2), .B(_13459__bF_buf3), .C(_13584_), .Y(_11355_) );
	INVX1 INVX1_1909 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .Y(_11356_) );
	NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_11356_), .B(_13458__bF_buf5), .C(_13466__bF_buf5), .Y(_11357_) );
	NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_13478__bF_buf1), .B(_11350_), .Y(_11358_) );
	OAI21X1 OAI21X1_4700 ( .gnd(gnd), .vdd(vdd), .A(_11351_), .B(_13478__bF_buf0), .C(_11358_), .Y(_11359_) );
	NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11359_), .C(_11355_), .Y(_11360_) );
	NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_11354_), .B(_11360_), .Y(_11361_) );
	INVX1 INVX1_1910 ( .gnd(gnd), .vdd(vdd), .A(_11298_), .Y(_11362_) );
	NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(_11313_), .B(_11319_), .C(_11314_), .Y(_11363_) );
	AOI21X1 AOI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_11362_), .B(_11363_), .C(_11320_), .Y(_11364_) );
	INVX1 INVX1_1911 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .Y(_11365_) );
	NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(_11363_), .B(_11365_), .C(_11301_), .Y(_11366_) );
	OAI21X1 OAI21X1_4701 ( .gnd(gnd), .vdd(vdd), .A(_11366_), .B(_13978_), .C(_11364_), .Y(_11367_) );
	XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_11367_), .B(_11361_), .Y(_11368_) );
	NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf3), .B(_11368_), .Y(_11369_) );
	NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_13584_), .B(_13687__bF_buf3), .Y(_11370_) );
	OAI21X1 OAI21X1_4702 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_10_), .B(_13687__bF_buf2), .C(_11370_), .Y(_11371_) );
	NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11355_), .Y(_11372_) );
	INVX1 INVX1_1912 ( .gnd(gnd), .vdd(vdd), .A(_11372_), .Y(_11373_) );
	OAI21X1 OAI21X1_4703 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf2), .B(csr_gpr_iu_ins_dec_xorp), .C(csr_gpr_iu_rs2_10_), .Y(_11374_) );
	OAI21X1 OAI21X1_4704 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(_13471_), .C(_11374_), .Y(_11375_) );
	OAI21X1 OAI21X1_4705 ( .gnd(gnd), .vdd(vdd), .A(_11375_), .B(_11373_), .C(amoxor_bF_buf1), .Y(_11376_) );
	AOI21X1 AOI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_11373_), .B(_11375_), .C(_11376_), .Y(_11377_) );
	OAI21X1 OAI21X1_4706 ( .gnd(gnd), .vdd(vdd), .A(_11351_), .B(_13776__bF_buf0), .C(_13454__bF_buf4), .Y(_11378_) );
	NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_11378_), .B(_11377_), .Y(_11379_) );
	OAI21X1 OAI21X1_4707 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf2), .B(_11371_), .C(_11379_), .Y(_11380_) );
	INVX1 INVX1_1913 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_10_), .Y(_11381_) );
	AOI21X1 AOI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_13397__bF_buf3), .C(_13398__bF_buf6), .Y(_11382_) );
	OAI21X1 OAI21X1_4708 ( .gnd(gnd), .vdd(vdd), .A(_11369_), .B(_11380_), .C(_11382_), .Y(_11383_) );
	NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_11351_), .B(_13695__bF_buf3), .Y(_11384_) );
	AOI21X1 AOI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_11384_), .B(_13694__bF_buf0), .C(_13391__bF_buf7), .Y(_11385_) );
	OAI21X1 OAI21X1_4709 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_10_), .B(_13392__bF_buf2), .C(_13412__bF_buf4), .Y(_11386_) );
	AOI21X1 AOI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_11383_), .B(_11385_), .C(_11386_), .Y(_11293__10_) );
	NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_11353_), .B(_11372_), .Y(_11387_) );
	AOI21X1 AOI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_11367_), .B(_11387_), .C(_11354_), .Y(_11388_) );
	OAI21X1 OAI21X1_4710 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf4), .C(_13589_), .Y(_11389_) );
	INVX1 INVX1_1914 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_11_), .Y(_11390_) );
	NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_11390_), .B(_13459__bF_buf1), .C(_13462__bF_buf1), .Y(_11391_) );
	NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(biu_pc_11_), .Y(_11392_) );
	INVX1 INVX1_1915 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .Y(_11393_) );
	OAI21X1 OAI21X1_4711 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(biu_ins_31_bF_buf2), .C(_13478__bF_buf4), .Y(_11394_) );
	OAI22X1 OAI22X1_819 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .B(_13478__bF_buf3), .C(_11392_), .D(_11394_), .Y(_11395_) );
	NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(_11389_), .B(_11395_), .C(_11391_), .Y(_11396_) );
	OAI21X1 OAI21X1_4712 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf3), .C(biu_biu_data_out_11_), .Y(_11397_) );
	NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_11_), .B(_13459__bF_buf0), .C(_13462__bF_buf0), .Y(_11398_) );
	INVX1 INVX1_1916 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .Y(_11399_) );
	NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11399_), .Y(_11400_) );
	INVX1 INVX1_1917 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .Y(_11401_) );
	AOI21X1 AOI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(_11401_), .C(_13707_), .Y(_11402_) );
	AOI22X1 AOI22X1_654 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_13707_), .C(_11400_), .D(_11402__bF_buf3), .Y(_11403_) );
	NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(_11397_), .B(_11403_), .C(_11398_), .Y(_11404_) );
	AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11404_), .Y(_11405_) );
	XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_11388_), .B(_11405_), .Y(_11406_) );
	AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_11406_), .B(_13489_), .Y(_11407_) );
	OAI21X1 OAI21X1_4713 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_13687__bF_buf1), .C(_13458__bF_buf2), .Y(_11408_) );
	AOI21X1 AOI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13687__bF_buf0), .C(_11408_), .Y(_11409_) );
	OAI21X1 OAI21X1_4714 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_11_), .B(_13476__bF_buf3), .C(_11391_), .Y(_11410_) );
	NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(_13471_), .Y(_11411_) );
	INVX4 INVX4_54 ( .gnd(gnd), .vdd(vdd), .A(_11411_), .Y(_11412_) );
	OAI21X1 OAI21X1_4715 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_13470__bF_buf2), .C(_11412__bF_buf3), .Y(_11413_) );
	AOI21X1 AOI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_11410_), .B(_11413_), .C(_13464__bF_buf3), .Y(_11414_) );
	OAI21X1 OAI21X1_4716 ( .gnd(gnd), .vdd(vdd), .A(_11410_), .B(_11413_), .C(_11414_), .Y(_11415_) );
	OAI21X1 OAI21X1_4717 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .B(_13776__bF_buf3), .C(_11415_), .Y(_11416_) );
	NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .B(_11409_), .Y(_11417_) );
	NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf3), .B(_11417_), .Y(_11418_) );
	INVX1 INVX1_1918 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_11_), .Y(_11419_) );
	AOI21X1 AOI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_11419_), .B(_13397__bF_buf2), .C(_13398__bF_buf5), .Y(_11420_) );
	OAI21X1 OAI21X1_4718 ( .gnd(gnd), .vdd(vdd), .A(_11407_), .B(_11418_), .C(_11420_), .Y(_11421_) );
	NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .B(_13695__bF_buf2), .Y(_11422_) );
	AOI21X1 AOI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_11422_), .B(_13694__bF_buf4), .C(_13391__bF_buf6), .Y(_11423_) );
	OAI21X1 OAI21X1_4719 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_11_), .B(_13392__bF_buf1), .C(_13412__bF_buf3), .Y(_11424_) );
	AOI21X1 AOI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_11421_), .B(_11423_), .C(_11424_), .Y(_11293__11_) );
	OAI21X1 OAI21X1_4720 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11355_), .C(_11359_), .Y(_11425_) );
	NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(_11425_), .B(_11387_), .C(_11405_), .Y(_11426_) );
	INVX1 INVX1_1919 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .Y(_11427_) );
	AOI21X1 AOI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_11354_), .B(_11404_), .C(_11427_), .Y(_11428_) );
	OAI21X1 OAI21X1_4721 ( .gnd(gnd), .vdd(vdd), .A(_11364_), .B(_11426_), .C(_11428_), .Y(_11429_) );
	NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11325_), .C(_11311_), .Y(_11430_) );
	NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11404_), .Y(_11431_) );
	NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_11354_), .B(_11360_), .C(_11431_), .Y(_11432_) );
	NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_11430_), .B(_11432_), .Y(_11433_) );
	NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_11433_), .B(_13978_), .Y(_11434_) );
	INVX1 INVX1_1920 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .Y(_11435_) );
	OAI21X1 OAI21X1_4722 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf2), .C(biu_biu_data_out_12_), .Y(_11436_) );
	OAI21X1 OAI21X1_4723 ( .gnd(gnd), .vdd(vdd), .A(_11435_), .B(_13463__bF_buf0), .C(_11436_), .Y(_11437_) );
	OAI21X1 OAI21X1_4724 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(biu_pc_12_), .C(_11402__bF_buf2), .Y(_11438_) );
	OAI21X1 OAI21X1_4725 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_13478__bF_buf2), .C(_11438_), .Y(_11439_) );
	NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_11439_), .B(_11437_), .Y(_11440_) );
	NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .B(_13476__bF_buf2), .Y(_11441_) );
	OAI21X1 OAI21X1_4726 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf0), .B(addp_bF_buf0), .C(csr_gpr_iu_rs2_12_), .Y(_11442_) );
	AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_11438_), .B(_11442_), .Y(_11443_) );
	NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .B(_11441_), .C(_11443_), .Y(_11444_) );
	AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(_11440_), .B(_11444_), .Y(_11445_) );
	OAI21X1 OAI21X1_4727 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11434_), .C(_11445_), .Y(_11446_) );
	NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11434_), .Y(_11447_) );
	NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_11444_), .B(_11440_), .Y(_11448_) );
	NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_11448_), .B(_11447_), .Y(_11449_) );
	NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_11446_), .B(_11449_), .Y(_11450_) );
	NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf2), .B(_11450_), .Y(_11451_) );
	NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_13580_), .B(_13687__bF_buf7), .Y(_11452_) );
	OAI21X1 OAI21X1_4728 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_13687__bF_buf6), .C(_11452_), .Y(_11453_) );
	AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_11441_), .B(_11436_), .Y(_11454_) );
	OAI21X1 OAI21X1_4729 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_13470__bF_buf1), .C(_11412__bF_buf2), .Y(_11455_) );
	OAI21X1 OAI21X1_4730 ( .gnd(gnd), .vdd(vdd), .A(_11455_), .B(_11454_), .C(amoxor_bF_buf0), .Y(_11456_) );
	AOI21X1 AOI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_11455_), .C(_11456_), .Y(_11457_) );
	OAI21X1 OAI21X1_4731 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_13776__bF_buf2), .C(_13454__bF_buf2), .Y(_11458_) );
	NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_11458_), .B(_11457_), .Y(_11459_) );
	OAI21X1 OAI21X1_4732 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf4), .B(_11453_), .C(_11459_), .Y(_11460_) );
	INVX1 INVX1_1921 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_12_), .Y(_11461_) );
	AOI21X1 AOI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_11461_), .B(_13397__bF_buf1), .C(_13398__bF_buf4), .Y(_11462_) );
	OAI21X1 OAI21X1_4733 ( .gnd(gnd), .vdd(vdd), .A(_11451_), .B(_11460_), .C(_11462_), .Y(_11463_) );
	NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_13695__bF_buf1), .Y(_11464_) );
	AOI21X1 AOI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_11464_), .B(_13694__bF_buf3), .C(_13391__bF_buf5), .Y(_11465_) );
	OAI21X1 OAI21X1_4734 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_12_), .B(_13392__bF_buf0), .C(_13412__bF_buf2), .Y(_11466_) );
	AOI21X1 AOI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_11463_), .B(_11465_), .C(_11466_), .Y(_11293__12_) );
	OAI21X1 OAI21X1_4735 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_11443_), .C(_11446_), .Y(_11467_) );
	OAI21X1 OAI21X1_4736 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf1), .C(_13563_), .Y(_11468_) );
	INVX1 INVX1_1922 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .Y(_11469_) );
	NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_11469_), .B(_13476__bF_buf1), .Y(_11470_) );
	INVX1 INVX1_1923 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .Y(_11471_) );
	NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11471_), .Y(_11472_) );
	AOI22X1 AOI22X1_655 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_13707_), .C(_11472_), .D(_11402__bF_buf1), .Y(_11473_) );
	INVX1 INVX1_1924 ( .gnd(gnd), .vdd(vdd), .A(_11473_), .Y(_11474_) );
	NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(_11468_), .B(_11470_), .C(_11474_), .Y(_11475_) );
	OAI21X1 OAI21X1_4737 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf8), .B(_13466__bF_buf0), .C(biu_biu_data_out_13_), .Y(_11476_) );
	NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .B(_13476__bF_buf0), .Y(_11477_) );
	NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(_11476_), .B(_11473_), .C(_11477_), .Y(_11478_) );
	AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_11475_), .B(_11478_), .Y(_11479_) );
	XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_11467_), .B(_11479_), .Y(_11480_) );
	NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf1), .B(_11480_), .Y(_11481_) );
	OAI21X1 OAI21X1_4738 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_13687__bF_buf5), .C(_13458__bF_buf7), .Y(_11482_) );
	AOI21X1 AOI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_13563_), .B(_13687__bF_buf4), .C(_11482_), .Y(_11483_) );
	OAI21X1 OAI21X1_4739 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .B(_13463__bF_buf4), .C(_11468_), .Y(_11484_) );
	OAI21X1 OAI21X1_4740 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_13470__bF_buf0), .C(_11412__bF_buf1), .Y(_11485_) );
	AOI21X1 AOI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_11484_), .B(_11485_), .C(_13464__bF_buf2), .Y(_11486_) );
	OAI21X1 OAI21X1_4741 ( .gnd(gnd), .vdd(vdd), .A(_11484_), .B(_11485_), .C(_11486_), .Y(_11487_) );
	OAI21X1 OAI21X1_4742 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_13776__bF_buf1), .C(_11487_), .Y(_11488_) );
	NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_11488_), .B(_11483_), .Y(_11489_) );
	NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf1), .B(_11489_), .Y(_11490_) );
	INVX1 INVX1_1925 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_13_), .Y(_11491_) );
	AOI21X1 AOI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_11491_), .B(_13397__bF_buf0), .C(_13398__bF_buf3), .Y(_11492_) );
	OAI21X1 OAI21X1_4743 ( .gnd(gnd), .vdd(vdd), .A(_11481_), .B(_11490_), .C(_11492_), .Y(_11493_) );
	NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_13695__bF_buf0), .Y(_11494_) );
	AOI21X1 AOI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_11494_), .B(_13694__bF_buf2), .C(_13391__bF_buf4), .Y(_11495_) );
	OAI21X1 OAI21X1_4744 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_13_), .B(_13392__bF_buf7), .C(_13412__bF_buf1), .Y(_11496_) );
	AOI21X1 AOI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_11493_), .B(_11495_), .C(_11496_), .Y(_11293__13_) );
	OAI21X1 OAI21X1_4745 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf6), .C(biu_biu_data_out_14_), .Y(_11497_) );
	NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_14_), .B(_13459__bF_buf3), .C(_13462__bF_buf3), .Y(_11498_) );
	INVX4 INVX4_55 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .Y(_11499_) );
	NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(biu_pc_14_), .Y(_11500_) );
	OAI22X1 OAI22X1_820 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_13478__bF_buf1), .C(_11500_), .D(_11394_), .Y(_11501_) );
	NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11501_), .C(_11498_), .Y(_11502_) );
	OAI21X1 OAI21X1_4746 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf5), .B(_13466__bF_buf5), .C(_13567_), .Y(_11503_) );
	INVX1 INVX1_1926 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_14_), .Y(_11504_) );
	NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(_11504_), .B(_13459__bF_buf2), .C(_13462__bF_buf2), .Y(_11505_) );
	INVX1 INVX1_1927 ( .gnd(gnd), .vdd(vdd), .A(_11500_), .Y(_11506_) );
	AOI22X1 AOI22X1_656 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_13707_), .C(_11506_), .D(_11402__bF_buf0), .Y(_11507_) );
	NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(_11503_), .B(_11507_), .C(_11505_), .Y(_11508_) );
	NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_11502_), .B(_11508_), .Y(_11509_) );
	AOI21X1 AOI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_11441_), .B(_11436_), .C(_11443_), .Y(_11510_) );
	INVX1 INVX1_1928 ( .gnd(gnd), .vdd(vdd), .A(_11475_), .Y(_11511_) );
	AOI21X1 AOI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_11510_), .B(_11478_), .C(_11511_), .Y(_11512_) );
	NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_11478_), .B(_11475_), .Y(_11513_) );
	NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_11513_), .B(_11448_), .Y(_11514_) );
	OAI21X1 OAI21X1_4747 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11434_), .C(_11514_), .Y(_11515_) );
	NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_11509_), .B(_11512_), .C(_11515_), .Y(_11516_) );
	INVX1 INVX1_1929 ( .gnd(gnd), .vdd(vdd), .A(_11509_), .Y(_11517_) );
	NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_11512_), .B(_11515_), .Y(_11518_) );
	NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_11517_), .B(_11518_), .Y(_11519_) );
	AOI21X1 AOI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_11519_), .B(_11516_), .C(_13488__bF_buf0), .Y(_11520_) );
	NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_14_), .B(_13687__bF_buf3), .Y(_11521_) );
	OAI21X1 OAI21X1_4748 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_13687__bF_buf2), .C(_11521_), .Y(_11522_) );
	OAI21X1 OAI21X1_4749 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_14_), .B(_13476__bF_buf3), .C(_11505_), .Y(_11523_) );
	OAI21X1 OAI21X1_4750 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_13470__bF_buf4), .C(_11412__bF_buf0), .Y(_11524_) );
	AOI21X1 AOI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_11523_), .B(_11524_), .C(_13464__bF_buf1), .Y(_11525_) );
	OAI21X1 OAI21X1_4751 ( .gnd(gnd), .vdd(vdd), .A(_11523_), .B(_11524_), .C(_11525_), .Y(_11526_) );
	OAI21X1 OAI21X1_4752 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_13776__bF_buf0), .C(_11526_), .Y(_11527_) );
	AOI21X1 AOI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_11522_), .B(_13458__bF_buf4), .C(_11527_), .Y(_11528_) );
	NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf0), .B(_11528_), .Y(_11529_) );
	INVX1 INVX1_1930 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_14_), .Y(_11530_) );
	AOI21X1 AOI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_11530_), .B(_13397__bF_buf4), .C(_13398__bF_buf2), .Y(_11531_) );
	OAI21X1 OAI21X1_4753 ( .gnd(gnd), .vdd(vdd), .A(_11520_), .B(_11529_), .C(_11531_), .Y(_11532_) );
	NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_13695__bF_buf5), .Y(_11533_) );
	AOI21X1 AOI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_11533_), .B(_13694__bF_buf1), .C(_13391__bF_buf3), .Y(_11534_) );
	OAI21X1 OAI21X1_4754 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_14_), .B(_13392__bF_buf6), .C(_13412__bF_buf0), .Y(_11535_) );
	AOI21X1 AOI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_11532_), .B(_11534_), .C(_11535_), .Y(_11293__14_) );
	NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11523_), .Y(_11536_) );
	AOI21X1 AOI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_11515_), .B(_11512_), .C(_11517_), .Y(_11537_) );
	NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11537_), .Y(_11538_) );
	OAI21X1 OAI21X1_4755 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf4), .C(_13572_), .Y(_11539_) );
	INVX1 INVX1_1931 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_15_), .Y(_11540_) );
	NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(_11540_), .B(_13459__bF_buf1), .C(_13462__bF_buf1), .Y(_11541_) );
	NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(biu_pc_15_), .Y(_11542_) );
	OAI22X1 OAI22X1_821 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13478__bF_buf0), .C(_11542_), .D(_11394_), .Y(_11543_) );
	NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(_11539_), .B(_11543_), .C(_11541_), .Y(_11544_) );
	OAI21X1 OAI21X1_4756 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf2), .B(_13466__bF_buf3), .C(biu_biu_data_out_15_), .Y(_11545_) );
	NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_15_), .B(_13459__bF_buf0), .C(_13462__bF_buf0), .Y(_11546_) );
	INVX1 INVX1_1932 ( .gnd(gnd), .vdd(vdd), .A(_11542_), .Y(_11547_) );
	AOI22X1 AOI22X1_657 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_13707_), .C(_11547_), .D(_11402__bF_buf3), .Y(_11548_) );
	NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(_11545_), .B(_11548_), .C(_11546_), .Y(_11549_) );
	NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(_11544_), .B(_11549_), .C(_11538_), .Y(_11550_) );
	NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_11544_), .B(_11549_), .Y(_11551_) );
	OAI21X1 OAI21X1_4757 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11537_), .C(_11551_), .Y(_11552_) );
	AOI21X1 AOI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_11550_), .B(_11552_), .C(_13488__bF_buf3), .Y(_11553_) );
	NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .B(_13687__bF_buf1), .Y(_11554_) );
	OAI21X1 OAI21X1_4758 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13687__bF_buf0), .C(_11554_), .Y(_11555_) );
	OAI21X1 OAI21X1_4759 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_15_), .B(_13476__bF_buf2), .C(_11541_), .Y(_11556_) );
	OAI21X1 OAI21X1_4760 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_13470__bF_buf3), .C(_11412__bF_buf3), .Y(_11557_) );
	AOI21X1 AOI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_11556_), .B(_11557_), .C(_13464__bF_buf0), .Y(_11558_) );
	OAI21X1 OAI21X1_4761 ( .gnd(gnd), .vdd(vdd), .A(_11556_), .B(_11557_), .C(_11558_), .Y(_11559_) );
	OAI21X1 OAI21X1_4762 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13776__bF_buf3), .C(_11559_), .Y(_11560_) );
	AOI21X1 AOI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_11555_), .B(_13458__bF_buf1), .C(_11560_), .Y(_11561_) );
	NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf4), .B(_11561_), .Y(_11562_) );
	INVX1 INVX1_1933 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_15_), .Y(_11563_) );
	AOI21X1 AOI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_11563_), .B(_13397__bF_buf3), .C(_13398__bF_buf1), .Y(_11564_) );
	OAI21X1 OAI21X1_4763 ( .gnd(gnd), .vdd(vdd), .A(_11553_), .B(_11562_), .C(_11564_), .Y(_11565_) );
	NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13695__bF_buf4), .Y(_11566_) );
	AOI21X1 AOI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_11566_), .B(_13694__bF_buf0), .C(_13391__bF_buf2), .Y(_11567_) );
	OAI21X1 OAI21X1_4764 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_15_), .B(_13392__bF_buf5), .C(_13412__bF_buf4), .Y(_11568_) );
	AOI21X1 AOI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_11565_), .B(_11567_), .C(_11568_), .Y(_11293__15_) );
	NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(_11544_), .B(_11549_), .C(_11509_), .Y(_11569_) );
	NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_11513_), .B(_11448_), .C(_11569_), .Y(_11570_) );
	NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_11430_), .B(_11432_), .C(_11570_), .Y(_11571_) );
	OAI21X1 OAI21X1_4765 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .B(_13476__bF_buf1), .C(_11546_), .Y(_11572_) );
	OAI21X1 OAI21X1_4766 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11523_), .C(_11544_), .Y(_11573_) );
	OAI21X1 OAI21X1_4767 ( .gnd(gnd), .vdd(vdd), .A(_11572_), .B(_11543_), .C(_11573_), .Y(_11574_) );
	OAI21X1 OAI21X1_4768 ( .gnd(gnd), .vdd(vdd), .A(_11569_), .B(_11512_), .C(_11574_), .Y(_11575_) );
	AOI21X1 AOI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11570_), .C(_11575_), .Y(_11576_) );
	OAI21X1 OAI21X1_4769 ( .gnd(gnd), .vdd(vdd), .A(_13978_), .B(_11571_), .C(_11576_), .Y(_11577_) );
	INVX1 INVX1_1934 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_16_), .Y(_11578_) );
	OAI21X1 OAI21X1_4770 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf2), .C(biu_biu_data_out_16_), .Y(_11579_) );
	OAI21X1 OAI21X1_4771 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_13463__bF_buf3), .C(_11579_), .Y(_11580_) );
	OAI21X1 OAI21X1_4772 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(biu_pc_16_), .C(_11402__bF_buf2), .Y(_11581_) );
	OAI21X1 OAI21X1_4773 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13478__bF_buf4), .C(_11581_), .Y(_11582_) );
	XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_11580_), .B(_11582_), .Y(_11583_) );
	XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_11577_), .B(_11583_), .Y(_11584_) );
	OAI21X1 OAI21X1_4774 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf3), .B(amoand), .C(_11584_), .Y(_11585_) );
	NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_16_), .B(_13687__bF_buf7), .Y(_11586_) );
	OAI21X1 OAI21X1_4775 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13687__bF_buf6), .C(_11586_), .Y(_11587_) );
	NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf8), .B(_11587_), .Y(_11588_) );
	MUX2X1 MUX2X1_168 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_16_), .B(biu_biu_data_out_16_), .S(_13476__bF_buf0), .Y(_11589_) );
	OAI21X1 OAI21X1_4776 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(_13470__bF_buf2), .C(_11412__bF_buf2), .Y(_11590_) );
	OAI21X1 OAI21X1_4777 ( .gnd(gnd), .vdd(vdd), .A(_11590_), .B(_11589_), .C(amoxor_bF_buf3), .Y(_11591_) );
	AOI21X1 AOI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_11589_), .B(_11590_), .C(_11591_), .Y(_11592_) );
	AOI21X1 AOI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(amoswap), .C(_11592_), .Y(_11593_) );
	NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(_11585_), .B(_11593_), .C(_11588_), .Y(_11594_) );
	INVX1 INVX1_1935 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_16_), .Y(_11595_) );
	AOI21X1 AOI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_11595_), .B(_13397__bF_buf2), .C(_13398__bF_buf0), .Y(_11596_) );
	OAI21X1 OAI21X1_4778 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_11594_), .C(_11596_), .Y(_11597_) );
	NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13695__bF_buf3), .Y(_11598_) );
	AOI21X1 AOI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_11598_), .B(_13694__bF_buf4), .C(_13391__bF_buf1), .Y(_11599_) );
	OAI21X1 OAI21X1_4779 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_16_), .B(_13392__bF_buf4), .C(_13412__bF_buf3), .Y(_11600_) );
	AOI21X1 AOI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_11597_), .B(_11599_), .C(_11600_), .Y(_11293__16_) );
	INVX1 INVX1_1936 ( .gnd(gnd), .vdd(vdd), .A(_11577_), .Y(_11601_) );
	NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_11582_), .B(_11580_), .Y(_11602_) );
	OAI21X1 OAI21X1_4780 ( .gnd(gnd), .vdd(vdd), .A(_11583_), .B(_11601_), .C(_11602_), .Y(_11603_) );
	INVX1 INVX1_1937 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_17_), .Y(_11604_) );
	OAI21X1 OAI21X1_4781 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf1), .C(biu_biu_data_out_17_), .Y(_11605_) );
	OAI21X1 OAI21X1_4782 ( .gnd(gnd), .vdd(vdd), .A(_11604_), .B(_13463__bF_buf2), .C(_11605_), .Y(_11606_) );
	INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .Y(_11607_) );
	OAI21X1 OAI21X1_4783 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(biu_pc_17_), .C(_11402__bF_buf1), .Y(_11608_) );
	OAI21X1 OAI21X1_4784 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_13478__bF_buf3), .C(_11608_), .Y(_11609_) );
	NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_11609_), .B(_11606_), .Y(_11610_) );
	OAI21X1 OAI21X1_4785 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf0), .C(_13553_), .Y(_11611_) );
	OAI21X1 OAI21X1_4786 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_17_), .B(_13463__bF_buf1), .C(_11611_), .Y(_11612_) );
	INVX1 INVX1_1938 ( .gnd(gnd), .vdd(vdd), .A(_11609_), .Y(_11613_) );
	NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_11612_), .B(_11613_), .Y(_11614_) );
	NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_11610_), .B(_11614_), .Y(_11615_) );
	XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11615_), .Y(_11616_) );
	AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_11616_), .B(_13489_), .Y(_11617_) );
	NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_17_), .B(_13687__bF_buf5), .Y(_11618_) );
	OAI21X1 OAI21X1_4787 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_13687__bF_buf4), .C(_11618_), .Y(_11619_) );
	OAI21X1 OAI21X1_4788 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_13470__bF_buf1), .C(_11412__bF_buf1), .Y(_11620_) );
	AOI21X1 AOI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_11612_), .B(_11620_), .C(_13464__bF_buf3), .Y(_11621_) );
	OAI21X1 OAI21X1_4789 ( .gnd(gnd), .vdd(vdd), .A(_11612_), .B(_11620_), .C(_11621_), .Y(_11622_) );
	OAI21X1 OAI21X1_4790 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_13776__bF_buf2), .C(_11622_), .Y(_11623_) );
	AOI21X1 AOI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_11619_), .B(_13458__bF_buf5), .C(_11623_), .Y(_11624_) );
	NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf3), .B(_11624_), .Y(_11625_) );
	INVX1 INVX1_1939 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_17_), .Y(_11626_) );
	AOI21X1 AOI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_11626_), .B(_13397__bF_buf1), .C(_13398__bF_buf6), .Y(_11627_) );
	OAI21X1 OAI21X1_4791 ( .gnd(gnd), .vdd(vdd), .A(_11617_), .B(_11625_), .C(_11627_), .Y(_11628_) );
	NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_13695__bF_buf2), .Y(_11629_) );
	AOI21X1 AOI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_11629_), .B(_13694__bF_buf3), .C(_13391__bF_buf0), .Y(_11630_) );
	OAI21X1 OAI21X1_4792 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_17_), .B(_13392__bF_buf3), .C(_13412__bF_buf2), .Y(_11631_) );
	AOI21X1 AOI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_11628_), .B(_11630_), .C(_11631_), .Y(_11293__17_) );
	OAI21X1 OAI21X1_4793 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf6), .C(_13543_), .Y(_11632_) );
	OAI21X1 OAI21X1_4794 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_18_), .B(_13463__bF_buf0), .C(_11632_), .Y(_11633_) );
	OAI21X1 OAI21X1_4795 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(biu_pc_18_), .C(_11402__bF_buf0), .Y(_11634_) );
	OAI21X1 OAI21X1_4796 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_13478__bF_buf2), .C(_11634_), .Y(_11635_) );
	NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_11635_), .B(_11633_), .Y(_11636_) );
	OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_11635_), .Y(_11637_) );
	NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .B(_11637_), .Y(_11638_) );
	OAI21X1 OAI21X1_4797 ( .gnd(gnd), .vdd(vdd), .A(_11602_), .B(_11615_), .C(_11610_), .Y(_11639_) );
	OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_11583_), .B(_11615_), .Y(_11640_) );
	NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_11640_), .B(_11601_), .Y(_11641_) );
	OAI21X1 OAI21X1_4798 ( .gnd(gnd), .vdd(vdd), .A(_11639_), .B(_11641_), .C(_11638_), .Y(_11642_) );
	INVX1 INVX1_1940 ( .gnd(gnd), .vdd(vdd), .A(_11638_), .Y(_11643_) );
	NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_11639_), .B(_11641_), .Y(_11644_) );
	NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_11643_), .B(_11644_), .Y(_11645_) );
	AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_11645_), .B(_11642_), .Y(_11646_) );
	AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_11646_), .B(_13489_), .Y(_11647_) );
	OAI21X1 OAI21X1_4799 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_13687__bF_buf3), .C(_13458__bF_buf3), .Y(_11648_) );
	AOI21X1 AOI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_13543_), .B(_13687__bF_buf2), .C(_11648_), .Y(_11649_) );
	OAI21X1 OAI21X1_4800 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_13470__bF_buf0), .C(_11412__bF_buf0), .Y(_11650_) );
	AOI21X1 AOI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_11650_), .C(_13464__bF_buf2), .Y(_11651_) );
	OAI21X1 OAI21X1_4801 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_11650_), .C(_11651_), .Y(_11652_) );
	OAI21X1 OAI21X1_4802 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_13776__bF_buf1), .C(_11652_), .Y(_11653_) );
	NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_11653_), .B(_11649_), .Y(_11654_) );
	NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf2), .B(_11654_), .Y(_11655_) );
	INVX1 INVX1_1941 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_18_), .Y(_11656_) );
	AOI21X1 AOI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_11656_), .B(_13397__bF_buf0), .C(_13398__bF_buf5), .Y(_11657_) );
	OAI21X1 OAI21X1_4803 ( .gnd(gnd), .vdd(vdd), .A(_11647_), .B(_11655_), .C(_11657_), .Y(_11658_) );
	NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_13695__bF_buf1), .Y(_11659_) );
	AOI21X1 AOI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_13694__bF_buf2), .C(_13391__bF_buf7), .Y(_11660_) );
	OAI21X1 OAI21X1_4804 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_18_), .B(_13392__bF_buf2), .C(_13412__bF_buf1), .Y(_11661_) );
	AOI21X1 AOI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_11658_), .B(_11660_), .C(_11661_), .Y(_11293__18_) );
	INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .Y(_11662_) );
	NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_11635_), .B(_11662_), .Y(_11663_) );
	OAI21X1 OAI21X1_4805 ( .gnd(gnd), .vdd(vdd), .A(_11643_), .B(_11644_), .C(_11663_), .Y(_11664_) );
	OAI21X1 OAI21X1_4806 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf2), .B(_13466__bF_buf5), .C(_13547_), .Y(_11665_) );
	OAI21X1 OAI21X1_4807 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_19_), .B(_13463__bF_buf4), .C(_11665_), .Y(_11666_) );
	INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .Y(_11667_) );
	NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11667_), .Y(_11668_) );
	AOI22X1 AOI22X1_658 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_13707_), .C(_11668_), .D(_11402__bF_buf3), .Y(_11669_) );
	OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_11666_), .B(_11669_), .Y(_11670_) );
	NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_11669_), .B(_11666_), .Y(_11671_) );
	AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_11670_), .B(_11671_), .Y(_11672_) );
	XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_11664_), .B(_11672_), .Y(_11673_) );
	NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf2), .B(_11673_), .Y(_11674_) );
	OAI21X1 OAI21X1_4808 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_13687__bF_buf1), .C(_13458__bF_buf1), .Y(_11675_) );
	AOI21X1 AOI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_13547_), .B(_13687__bF_buf0), .C(_11675_), .Y(_11676_) );
	OAI21X1 OAI21X1_4809 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_13470__bF_buf4), .C(_11412__bF_buf3), .Y(_11677_) );
	AOI21X1 AOI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_11666_), .B(_11677_), .C(_13464__bF_buf1), .Y(_11678_) );
	OAI21X1 OAI21X1_4810 ( .gnd(gnd), .vdd(vdd), .A(_11666_), .B(_11677_), .C(_11678_), .Y(_11679_) );
	OAI21X1 OAI21X1_4811 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_13776__bF_buf0), .C(_11679_), .Y(_11680_) );
	NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_11680_), .B(_11676_), .Y(_11681_) );
	NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf1), .B(_11681_), .Y(_11682_) );
	INVX1 INVX1_1942 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_19_), .Y(_11683_) );
	AOI21X1 AOI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_11683_), .B(_13397__bF_buf4), .C(_13398__bF_buf4), .Y(_11684_) );
	OAI21X1 OAI21X1_4812 ( .gnd(gnd), .vdd(vdd), .A(_11674_), .B(_11682_), .C(_11684_), .Y(_11685_) );
	NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_13695__bF_buf0), .Y(_11686_) );
	AOI21X1 AOI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_11686_), .B(_13694__bF_buf1), .C(_13391__bF_buf6), .Y(_11687_) );
	OAI21X1 OAI21X1_4813 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_19_), .B(_13392__bF_buf1), .C(_13412__bF_buf0), .Y(_11688_) );
	AOI21X1 AOI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_11685_), .B(_11687_), .C(_11688_), .Y(_11293__19_) );
	NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_11671_), .B(_11670_), .Y(_11689_) );
	OAI21X1 OAI21X1_4814 ( .gnd(gnd), .vdd(vdd), .A(_11663_), .B(_11689_), .C(_11670_), .Y(_11690_) );
	AOI21X1 AOI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .B(_11637_), .C(_11689_), .Y(_11691_) );
	AOI21X1 AOI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_11691_), .B(_11639_), .C(_11690_), .Y(_11692_) );
	NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_11615_), .B(_11583_), .Y(_11693_) );
	NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_11693_), .B(_11691_), .Y(_11694_) );
	OAI21X1 OAI21X1_4815 ( .gnd(gnd), .vdd(vdd), .A(_11694_), .B(_11601_), .C(_11692_), .Y(_11695_) );
	INVX1 INVX1_1943 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_20_), .Y(_11696_) );
	OAI21X1 OAI21X1_4816 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf4), .C(biu_biu_data_out_20_), .Y(_11697_) );
	OAI21X1 OAI21X1_4817 ( .gnd(gnd), .vdd(vdd), .A(_11696_), .B(_13463__bF_buf3), .C(_11697_), .Y(_11698_) );
	INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .Y(_11699_) );
	OAI21X1 OAI21X1_4818 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(biu_pc_20_), .C(_11402__bF_buf2), .Y(_11700_) );
	OAI21X1 OAI21X1_4819 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_13478__bF_buf1), .C(_11700_), .Y(_11701_) );
	NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_11701_), .B(_11699_), .Y(_11702_) );
	INVX1 INVX1_1944 ( .gnd(gnd), .vdd(vdd), .A(_11701_), .Y(_11703_) );
	NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .B(_11703_), .Y(_11704_) );
	NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_11704_), .B(_11702_), .Y(_11705_) );
	XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_11695_), .B(_11705_), .Y(_11706_) );
	AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_11706_), .B(_13489_), .Y(_11707_) );
	NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_20_), .B(_13687__bF_buf7), .Y(_11708_) );
	OAI21X1 OAI21X1_4820 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_13687__bF_buf6), .C(_11708_), .Y(_11709_) );
	OAI21X1 OAI21X1_4821 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(_13470__bF_buf3), .C(_11412__bF_buf2), .Y(_11710_) );
	AOI21X1 AOI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11710_), .C(_13464__bF_buf0), .Y(_11711_) );
	OAI21X1 OAI21X1_4822 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11710_), .C(_11711_), .Y(_11712_) );
	OAI21X1 OAI21X1_4823 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_13776__bF_buf3), .C(_11712_), .Y(_11713_) );
	AOI21X1 AOI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_11709_), .B(_13458__bF_buf8), .C(_11713_), .Y(_11714_) );
	NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf0), .B(_11714_), .Y(_11715_) );
	INVX1 INVX1_1945 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_20_), .Y(_11716_) );
	AOI21X1 AOI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_11716_), .B(_13397__bF_buf3), .C(_13398__bF_buf3), .Y(_11717_) );
	OAI21X1 OAI21X1_4824 ( .gnd(gnd), .vdd(vdd), .A(_11707_), .B(_11715_), .C(_11717_), .Y(_11718_) );
	NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_13695__bF_buf5), .Y(_11719_) );
	AOI21X1 AOI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_11719_), .B(_13694__bF_buf0), .C(_13391__bF_buf5), .Y(_11720_) );
	OAI21X1 OAI21X1_4825 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_20_), .B(_13392__bF_buf0), .C(_13412__bF_buf4), .Y(_11721_) );
	AOI21X1 AOI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_11718_), .B(_11720_), .C(_11721_), .Y(_11293__20_) );
	NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_11705_), .B(_11695_), .Y(_11722_) );
	OAI21X1 OAI21X1_4826 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11703_), .C(_11722_), .Y(_11723_) );
	INVX1 INVX1_1946 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_21_), .Y(_11724_) );
	OAI21X1 OAI21X1_4827 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf3), .C(biu_biu_data_out_21_), .Y(_11725_) );
	OAI21X1 OAI21X1_4828 ( .gnd(gnd), .vdd(vdd), .A(_11724_), .B(_13463__bF_buf2), .C(_11725_), .Y(_11726_) );
	INVX4 INVX4_56 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .Y(_11727_) );
	OAI21X1 OAI21X1_4829 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(biu_pc_21_), .C(_11402__bF_buf1), .Y(_11728_) );
	OAI21X1 OAI21X1_4830 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_13478__bF_buf0), .C(_11728_), .Y(_11729_) );
	NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_11729_), .B(_11726_), .Y(_11730_) );
	OAI21X1 OAI21X1_4831 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf2), .C(_13523_), .Y(_11731_) );
	OAI21X1 OAI21X1_4832 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_21_), .B(_13463__bF_buf1), .C(_11731_), .Y(_11732_) );
	INVX1 INVX1_1947 ( .gnd(gnd), .vdd(vdd), .A(_11729_), .Y(_11733_) );
	NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11733_), .Y(_11734_) );
	NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_11730_), .B(_11734_), .Y(_11735_) );
	XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_11723_), .B(_11735_), .Y(_11736_) );
	AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_11736_), .B(_13489_), .Y(_11737_) );
	NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_21_), .B(_13687__bF_buf5), .Y(_11738_) );
	OAI21X1 OAI21X1_4833 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_13687__bF_buf4), .C(_11738_), .Y(_11739_) );
	OAI21X1 OAI21X1_4834 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_13470__bF_buf2), .C(_11412__bF_buf1), .Y(_11740_) );
	AOI21X1 AOI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11740_), .C(_13464__bF_buf3), .Y(_11741_) );
	OAI21X1 OAI21X1_4835 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11740_), .C(_11741_), .Y(_11742_) );
	OAI21X1 OAI21X1_4836 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_13776__bF_buf2), .C(_11742_), .Y(_11743_) );
	AOI21X1 AOI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_11739_), .B(_13458__bF_buf5), .C(_11743_), .Y(_11744_) );
	NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf4), .B(_11744_), .Y(_11745_) );
	INVX1 INVX1_1948 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_21_), .Y(_11746_) );
	AOI21X1 AOI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_11746_), .B(_13397__bF_buf2), .C(_13398__bF_buf2), .Y(_11747_) );
	OAI21X1 OAI21X1_4837 ( .gnd(gnd), .vdd(vdd), .A(_11737_), .B(_11745_), .C(_11747_), .Y(_11748_) );
	NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_13695__bF_buf4), .Y(_11749_) );
	AOI21X1 AOI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_11749_), .B(_13694__bF_buf4), .C(_13391__bF_buf4), .Y(_11750_) );
	OAI21X1 OAI21X1_4838 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_21_), .B(_13392__bF_buf7), .C(_13412__bF_buf3), .Y(_11751_) );
	AOI21X1 AOI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_11748_), .B(_11750_), .C(_11751_), .Y(_11293__21_) );
	OAI21X1 OAI21X1_4839 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf1), .C(_13531_), .Y(_11752_) );
	OAI21X1 OAI21X1_4840 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_22_), .B(_13463__bF_buf0), .C(_11752_), .Y(_11753_) );
	OAI21X1 OAI21X1_4841 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(biu_pc_22_), .C(_11402__bF_buf0), .Y(_11754_) );
	OAI21X1 OAI21X1_4842 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .B(_13478__bF_buf4), .C(_11754_), .Y(_11755_) );
	NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_11755_), .B(_11753_), .Y(_11756_) );
	INVX1 INVX1_1949 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_22_), .Y(_11757_) );
	OAI21X1 OAI21X1_4843 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf0), .C(biu_biu_data_out_22_), .Y(_11758_) );
	OAI21X1 OAI21X1_4844 ( .gnd(gnd), .vdd(vdd), .A(_11757_), .B(_13463__bF_buf4), .C(_11758_), .Y(_11759_) );
	OAI21X1 OAI21X1_4845 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf2), .B(addp_bF_buf4), .C(csr_gpr_iu_rs2_22_), .Y(_11760_) );
	AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_11754_), .B(_11760_), .Y(_11761_) );
	NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11759_), .Y(_11762_) );
	NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_11756_), .B(_11762_), .Y(_11763_) );
	NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_11701_), .B(_11698_), .Y(_11764_) );
	NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(_11764_), .B(_11730_), .C(_11722_), .Y(_11765_) );
	OAI21X1 OAI21X1_4846 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_11729_), .C(_11765_), .Y(_11766_) );
	NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .B(_11766_), .Y(_11767_) );
	OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_11766_), .B(_11763_), .Y(_11768_) );
	AOI21X1 AOI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_11768_), .B(_11767_), .C(_13488__bF_buf1), .Y(_11769_) );
	OAI21X1 OAI21X1_4847 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_13687__bF_buf3), .C(_13458__bF_buf2), .Y(_11770_) );
	AOI21X1 AOI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_13531_), .B(_13687__bF_buf2), .C(_11770_), .Y(_11771_) );
	OAI21X1 OAI21X1_4848 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_13470__bF_buf1), .C(_11412__bF_buf0), .Y(_11772_) );
	AOI21X1 AOI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_11753_), .B(_11772_), .C(_13464__bF_buf2), .Y(_11773_) );
	OAI21X1 OAI21X1_4849 ( .gnd(gnd), .vdd(vdd), .A(_11753_), .B(_11772_), .C(_11773_), .Y(_11774_) );
	OAI21X1 OAI21X1_4850 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .B(_13776__bF_buf1), .C(_11774_), .Y(_11775_) );
	NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .B(_11771_), .Y(_11776_) );
	NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf3), .B(_11776_), .Y(_11777_) );
	INVX1 INVX1_1950 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_22_), .Y(_11778_) );
	AOI21X1 AOI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_11778_), .B(_13397__bF_buf1), .C(_13398__bF_buf1), .Y(_11779_) );
	OAI21X1 OAI21X1_4851 ( .gnd(gnd), .vdd(vdd), .A(_11777_), .B(_11769_), .C(_11779_), .Y(_11780_) );
	NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .B(_13695__bF_buf3), .Y(_11781_) );
	AOI21X1 AOI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_11781_), .B(_13694__bF_buf3), .C(_13391__bF_buf3), .Y(_11782_) );
	OAI21X1 OAI21X1_4852 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_22_), .B(_13392__bF_buf6), .C(_13412__bF_buf2), .Y(_11783_) );
	AOI21X1 AOI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_11780_), .B(_11782_), .C(_11783_), .Y(_11293__22_) );
	NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11753_), .Y(_11784_) );
	INVX1 INVX1_1951 ( .gnd(gnd), .vdd(vdd), .A(_11784_), .Y(_11785_) );
	AOI21X1 AOI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_11702_), .B(_11704_), .C(_11735_), .Y(_11786_) );
	NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .B(_11695_), .Y(_11787_) );
	OAI21X1 OAI21X1_4853 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11733_), .C(_11764_), .Y(_11788_) );
	OAI21X1 OAI21X1_4854 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_11729_), .C(_11788_), .Y(_11789_) );
	AOI22X1 AOI22X1_659 ( .gnd(gnd), .vdd(vdd), .A(_11756_), .B(_11762_), .C(_11789_), .D(_11787_), .Y(_11790_) );
	INVX1 INVX1_1952 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .Y(_11791_) );
	OAI21X1 OAI21X1_4855 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf6), .C(_13528_), .Y(_11792_) );
	OAI21X1 OAI21X1_4856 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_23_), .B(_13463__bF_buf3), .C(_11792_), .Y(_11793_) );
	OAI21X1 OAI21X1_4857 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(biu_pc_23_), .C(_11402__bF_buf3), .Y(_11794_) );
	OAI21X1 OAI21X1_4858 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13478__bF_buf3), .C(_11794_), .Y(_11795_) );
	NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_11795_), .B(_11793_), .Y(_11796_) );
	INVX1 INVX1_1953 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_23_), .Y(_11797_) );
	OAI21X1 OAI21X1_4859 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf5), .C(biu_biu_data_out_23_), .Y(_11798_) );
	OAI21X1 OAI21X1_4860 ( .gnd(gnd), .vdd(vdd), .A(_11797_), .B(_13463__bF_buf2), .C(_11798_), .Y(_11799_) );
	OAI21X1 OAI21X1_4861 ( .gnd(gnd), .vdd(vdd), .A(amoadd_bF_buf1), .B(addp_bF_buf3), .C(csr_gpr_iu_rs2_23_), .Y(_11800_) );
	AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_11794_), .B(_11800_), .Y(_11801_) );
	NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_11801_), .B(_11799_), .Y(_11802_) );
	AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_11796_), .B(_11802_), .Y(_11803_) );
	NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(_11785_), .B(_11803_), .C(_11791_), .Y(_11804_) );
	NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_11796_), .B(_11802_), .Y(_11805_) );
	OAI21X1 OAI21X1_4862 ( .gnd(gnd), .vdd(vdd), .A(_11784_), .B(_11790_), .C(_11805_), .Y(_11806_) );
	NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_11806_), .B(_11804_), .Y(_11807_) );
	NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf0), .B(_11807_), .Y(_11808_) );
	NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_23_), .B(_13687__bF_buf1), .Y(_11809_) );
	OAI21X1 OAI21X1_4863 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13687__bF_buf0), .C(_11809_), .Y(_11810_) );
	OAI21X1 OAI21X1_4864 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_23_), .B(_13470__bF_buf0), .C(_11412__bF_buf3), .Y(_11811_) );
	AOI21X1 AOI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11811_), .C(_13464__bF_buf1), .Y(_11812_) );
	OAI21X1 OAI21X1_4865 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11811_), .C(_11812_), .Y(_11813_) );
	OAI21X1 OAI21X1_4866 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13776__bF_buf0), .C(_11813_), .Y(_11814_) );
	AOI21X1 AOI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_11810_), .B(_13458__bF_buf8), .C(_11814_), .Y(_11815_) );
	NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf2), .B(_11815_), .Y(_11816_) );
	INVX1 INVX1_1954 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_23_), .Y(_11817_) );
	AOI21X1 AOI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_11817_), .B(_13397__bF_buf0), .C(_13398__bF_buf0), .Y(_11818_) );
	OAI21X1 OAI21X1_4867 ( .gnd(gnd), .vdd(vdd), .A(_11816_), .B(_11808_), .C(_11818_), .Y(_11819_) );
	NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13695__bF_buf2), .Y(_11820_) );
	AOI21X1 AOI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_11820_), .B(_13694__bF_buf2), .C(_13391__bF_buf2), .Y(_11821_) );
	OAI21X1 OAI21X1_4868 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_23_), .B(_13392__bF_buf5), .C(_13412__bF_buf1), .Y(_11822_) );
	AOI21X1 AOI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_11819_), .B(_11821_), .C(_11822_), .Y(_11293__23_) );
	AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .B(_11805_), .Y(_11823_) );
	NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .B(_11823_), .Y(_11824_) );
	NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(_11694_), .Y(_11825_) );
	OAI21X1 OAI21X1_4869 ( .gnd(gnd), .vdd(vdd), .A(_11764_), .B(_11735_), .C(_11730_), .Y(_11826_) );
	NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_11795_), .B(_11799_), .Y(_11827_) );
	OAI21X1 OAI21X1_4870 ( .gnd(gnd), .vdd(vdd), .A(_11785_), .B(_11803_), .C(_11827_), .Y(_11828_) );
	AOI21X1 AOI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_11826_), .B(_11823_), .C(_11828_), .Y(_11829_) );
	OAI21X1 OAI21X1_4871 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(_11692_), .C(_11829_), .Y(_11830_) );
	AOI21X1 AOI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_11577_), .B(_11825_), .C(_11830_), .Y(_11831_) );
	INVX1 INVX1_1955 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_24_), .Y(_11832_) );
	OAI21X1 OAI21X1_4872 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf7), .B(_13466__bF_buf4), .C(biu_biu_data_out_24_), .Y(_11833_) );
	OAI21X1 OAI21X1_4873 ( .gnd(gnd), .vdd(vdd), .A(_11832_), .B(_13463__bF_buf1), .C(_11833_), .Y(_11834_) );
	OAI21X1 OAI21X1_4874 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(biu_pc_24_), .C(_11402__bF_buf2), .Y(_11835_) );
	OAI21X1 OAI21X1_4875 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13478__bF_buf2), .C(_11835_), .Y(_11836_) );
	XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(_11836_), .Y(_11837_) );
	XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_11831_), .B(_11837_), .Y(_11838_) );
	AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .B(_13489_), .Y(_11839_) );
	NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_24_), .B(_13687__bF_buf7), .Y(_11840_) );
	OAI21X1 OAI21X1_4876 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13687__bF_buf6), .C(_11840_), .Y(_11841_) );
	INVX1 INVX1_1956 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .Y(_11842_) );
	OAI21X1 OAI21X1_4877 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .B(_13470__bF_buf4), .C(_11412__bF_buf2), .Y(_11843_) );
	AOI21X1 AOI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_11842_), .B(_11843_), .C(_13464__bF_buf0), .Y(_11844_) );
	OAI21X1 OAI21X1_4878 ( .gnd(gnd), .vdd(vdd), .A(_11842_), .B(_11843_), .C(_11844_), .Y(_11845_) );
	OAI21X1 OAI21X1_4879 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13776__bF_buf3), .C(_11845_), .Y(_11846_) );
	AOI21X1 AOI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_11841_), .B(_13458__bF_buf6), .C(_11846_), .Y(_11847_) );
	NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf1), .B(_11847_), .Y(_11848_) );
	INVX1 INVX1_1957 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_24_), .Y(_11849_) );
	AOI21X1 AOI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .B(_13397__bF_buf4), .C(_13398__bF_buf6), .Y(_11850_) );
	OAI21X1 OAI21X1_4880 ( .gnd(gnd), .vdd(vdd), .A(_11839_), .B(_11848_), .C(_11850_), .Y(_11851_) );
	NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13695__bF_buf1), .Y(_11852_) );
	AOI21X1 AOI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .B(_13694__bF_buf1), .C(_13391__bF_buf1), .Y(_11853_) );
	OAI21X1 OAI21X1_4881 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_24_), .B(_13392__bF_buf4), .C(_13412__bF_buf0), .Y(_11854_) );
	AOI21X1 AOI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_11851_), .B(_11853_), .C(_11854_), .Y(_11293__24_) );
	NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_11836_), .B(_11834_), .Y(_11855_) );
	INVX1 INVX1_1958 ( .gnd(gnd), .vdd(vdd), .A(_11837_), .Y(_11856_) );
	OAI21X1 OAI21X1_4882 ( .gnd(gnd), .vdd(vdd), .A(_11856_), .B(_11831_), .C(_11855_), .Y(_11857_) );
	INVX1 INVX1_1959 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_25_), .Y(_11858_) );
	OAI21X1 OAI21X1_4883 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf5), .B(_13466__bF_buf3), .C(biu_biu_data_out_25_), .Y(_11859_) );
	OAI21X1 OAI21X1_4884 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_13463__bF_buf0), .C(_11859_), .Y(_11860_) );
	OAI21X1 OAI21X1_4885 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(biu_pc_25_), .C(_11402__bF_buf1), .Y(_11861_) );
	OAI21X1 OAI21X1_4886 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_13478__bF_buf1), .C(_11861_), .Y(_11862_) );
	NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_11862_), .B(_11860_), .Y(_11863_) );
	INVX1 INVX1_1960 ( .gnd(gnd), .vdd(vdd), .A(_11863_), .Y(_11864_) );
	NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_11862_), .B(_11860_), .Y(_11865_) );
	NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_11865_), .B(_11864_), .Y(_11866_) );
	XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11866_), .Y(_11867_) );
	NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf3), .B(_11867_), .Y(_11868_) );
	NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_25_), .B(_13687__bF_buf5), .Y(_11869_) );
	OAI21X1 OAI21X1_4887 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_13687__bF_buf4), .C(_11869_), .Y(_11870_) );
	INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .Y(_11871_) );
	OAI21X1 OAI21X1_4888 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_13470__bF_buf3), .C(_11412__bF_buf1), .Y(_11872_) );
	AOI21X1 AOI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_11871_), .B(_11872_), .C(_13464__bF_buf3), .Y(_11873_) );
	OAI21X1 OAI21X1_4889 ( .gnd(gnd), .vdd(vdd), .A(_11871_), .B(_11872_), .C(_11873_), .Y(_11874_) );
	OAI21X1 OAI21X1_4890 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_13776__bF_buf2), .C(_11874_), .Y(_11875_) );
	AOI21X1 AOI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_11870_), .B(_13458__bF_buf4), .C(_11875_), .Y(_11876_) );
	NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf0), .B(_11876_), .Y(_11877_) );
	INVX1 INVX1_1961 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_25_), .Y(_11878_) );
	AOI21X1 AOI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_11878_), .B(_13397__bF_buf3), .C(_13398__bF_buf5), .Y(_11879_) );
	OAI21X1 OAI21X1_4891 ( .gnd(gnd), .vdd(vdd), .A(_11868_), .B(_11877_), .C(_11879_), .Y(_11880_) );
	NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_13695__bF_buf0), .Y(_11881_) );
	AOI21X1 AOI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_11881_), .B(_13694__bF_buf0), .C(_13391__bF_buf0), .Y(_11882_) );
	OAI21X1 OAI21X1_4892 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_25_), .B(_13392__bF_buf3), .C(_13412__bF_buf4), .Y(_11883_) );
	AOI21X1 AOI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_11880_), .B(_11882_), .C(_11883_), .Y(_11293__25_) );
	INVX1 INVX1_1962 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_26_), .Y(_11884_) );
	OAI21X1 OAI21X1_4893 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf3), .B(_13466__bF_buf2), .C(biu_biu_data_out_26_), .Y(_11885_) );
	OAI21X1 OAI21X1_4894 ( .gnd(gnd), .vdd(vdd), .A(_11884_), .B(_13463__bF_buf4), .C(_11885_), .Y(_11886_) );
	INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .Y(_11887_) );
	OAI21X1 OAI21X1_4895 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(biu_pc_26_), .C(_11402__bF_buf0), .Y(_11888_) );
	OAI21X1 OAI21X1_4896 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_13478__bF_buf0), .C(_11888_), .Y(_11889_) );
	NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .B(_11886_), .Y(_11890_) );
	INVX1 INVX1_1963 ( .gnd(gnd), .vdd(vdd), .A(_11890_), .Y(_11891_) );
	NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .B(_11886_), .Y(_11892_) );
	NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_11892_), .B(_11891_), .Y(_11893_) );
	OAI21X1 OAI21X1_4897 ( .gnd(gnd), .vdd(vdd), .A(_11855_), .B(_11865_), .C(_11863_), .Y(_11894_) );
	NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_11837_), .B(_11866_), .Y(_11895_) );
	NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_11895_), .B(_11831_), .Y(_11896_) );
	OAI21X1 OAI21X1_4898 ( .gnd(gnd), .vdd(vdd), .A(_11894_), .B(_11896_), .C(_11893_), .Y(_11897_) );
	NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_11894_), .B(_11896_), .Y(_11898_) );
	OAI21X1 OAI21X1_4899 ( .gnd(gnd), .vdd(vdd), .A(_11891_), .B(_11892_), .C(_11898_), .Y(_11899_) );
	NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_11897_), .B(_11899_), .Y(_11900_) );
	NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf2), .B(_11900_), .Y(_11901_) );
	OAI21X1 OAI21X1_4900 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_13687__bF_buf3), .C(_13458__bF_buf2), .Y(_11902_) );
	AOI21X1 AOI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_13507_), .B(_13687__bF_buf2), .C(_11902_), .Y(_11903_) );
	INVX1 INVX1_1964 ( .gnd(gnd), .vdd(vdd), .A(_11886_), .Y(_11904_) );
	OAI21X1 OAI21X1_4901 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_13470__bF_buf2), .C(_11412__bF_buf0), .Y(_11905_) );
	AOI21X1 AOI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_11904_), .B(_11905_), .C(_13464__bF_buf2), .Y(_11906_) );
	OAI21X1 OAI21X1_4902 ( .gnd(gnd), .vdd(vdd), .A(_11904_), .B(_11905_), .C(_11906_), .Y(_11907_) );
	OAI21X1 OAI21X1_4903 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_13776__bF_buf1), .C(_11907_), .Y(_11908_) );
	NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_11908_), .B(_11903_), .Y(_11909_) );
	NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf4), .B(_11909_), .Y(_11910_) );
	INVX1 INVX1_1965 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_26_), .Y(_11911_) );
	AOI21X1 AOI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_11911_), .B(_13397__bF_buf2), .C(_13398__bF_buf4), .Y(_11912_) );
	OAI21X1 OAI21X1_4904 ( .gnd(gnd), .vdd(vdd), .A(_11901_), .B(_11910_), .C(_11912_), .Y(_11913_) );
	NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_13695__bF_buf5), .Y(_11914_) );
	AOI21X1 AOI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_11914_), .B(_13694__bF_buf4), .C(_13391__bF_buf7), .Y(_11915_) );
	OAI21X1 OAI21X1_4905 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_26_), .B(_13392__bF_buf2), .C(_13412__bF_buf3), .Y(_11916_) );
	AOI21X1 AOI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_11913_), .B(_11915_), .C(_11916_), .Y(_11293__26_) );
	INVX1 INVX1_1966 ( .gnd(gnd), .vdd(vdd), .A(_11893_), .Y(_11917_) );
	OAI21X1 OAI21X1_4906 ( .gnd(gnd), .vdd(vdd), .A(_11917_), .B(_11898_), .C(_11890_), .Y(_11918_) );
	INVX1 INVX1_1967 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_27_), .Y(_11919_) );
	OAI21X1 OAI21X1_4907 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf1), .C(biu_biu_data_out_27_), .Y(_11920_) );
	OAI21X1 OAI21X1_4908 ( .gnd(gnd), .vdd(vdd), .A(_11919_), .B(_13463__bF_buf3), .C(_11920_), .Y(_11921_) );
	OAI21X1 OAI21X1_4909 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(biu_pc_27_), .C(_11402__bF_buf3), .Y(_11922_) );
	OAI21X1 OAI21X1_4910 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13478__bF_buf4), .C(_11922_), .Y(_11923_) );
	NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_11923_), .B(_11921_), .Y(_11924_) );
	OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .B(_11923_), .Y(_11925_) );
	NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_11924_), .B(_11925_), .Y(_11926_) );
	OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_11918_), .B(_11926_), .Y(_11927_) );
	NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_11918_), .Y(_11928_) );
	AOI21X1 AOI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_11927_), .B(_11928_), .C(_13488__bF_buf1), .Y(_11929_) );
	NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_27_), .B(_13687__bF_buf1), .Y(_11930_) );
	OAI21X1 OAI21X1_4911 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13687__bF_buf0), .C(_11930_), .Y(_11931_) );
	INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .Y(_11932_) );
	OAI21X1 OAI21X1_4912 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_27_), .B(_13470__bF_buf1), .C(_11412__bF_buf3), .Y(_11933_) );
	AOI21X1 AOI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_11933_), .C(_13464__bF_buf1), .Y(_11934_) );
	OAI21X1 OAI21X1_4913 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_11933_), .C(_11934_), .Y(_11935_) );
	OAI21X1 OAI21X1_4914 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13776__bF_buf0), .C(_11935_), .Y(_11936_) );
	AOI21X1 AOI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_11931_), .B(_13458__bF_buf0), .C(_11936_), .Y(_11937_) );
	NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf3), .B(_11937_), .Y(_11938_) );
	INVX1 INVX1_1968 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_27_), .Y(_11939_) );
	AOI21X1 AOI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_13397__bF_buf1), .C(_13398__bF_buf3), .Y(_11940_) );
	OAI21X1 OAI21X1_4915 ( .gnd(gnd), .vdd(vdd), .A(_11938_), .B(_11929_), .C(_11940_), .Y(_11941_) );
	NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13695__bF_buf4), .Y(_11942_) );
	AOI21X1 AOI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_11942_), .B(_13694__bF_buf3), .C(_13391__bF_buf6), .Y(_11943_) );
	OAI21X1 OAI21X1_4916 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_27_), .B(_13392__bF_buf1), .C(_13412__bF_buf2), .Y(_11944_) );
	AOI21X1 AOI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_11941_), .B(_11943_), .C(_11944_), .Y(_11293__27_) );
	NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_11917_), .Y(_11945_) );
	INVX1 INVX1_1969 ( .gnd(gnd), .vdd(vdd), .A(_11945_), .Y(_11946_) );
	OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_11946_), .B(_11895_), .Y(_11947_) );
	OAI21X1 OAI21X1_4917 ( .gnd(gnd), .vdd(vdd), .A(_11890_), .B(_11926_), .C(_11924_), .Y(_11948_) );
	AOI21X1 AOI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_11945_), .B(_11894_), .C(_11948_), .Y(_11949_) );
	OAI21X1 OAI21X1_4918 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .B(_11831_), .C(_11949_), .Y(_11950_) );
	INVX1 INVX1_1970 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_28_), .Y(_11951_) );
	OAI21X1 OAI21X1_4919 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf8), .B(_13466__bF_buf0), .C(biu_biu_data_out_28_), .Y(_11952_) );
	OAI21X1 OAI21X1_4920 ( .gnd(gnd), .vdd(vdd), .A(_11951_), .B(_13463__bF_buf2), .C(_11952_), .Y(_11953_) );
	INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .Y(_11954_) );
	INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .Y(_11955_) );
	OAI21X1 OAI21X1_4921 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(biu_pc_28_), .C(_11402__bF_buf2), .Y(_11956_) );
	OAI21X1 OAI21X1_4922 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_13478__bF_buf3), .C(_11956_), .Y(_11957_) );
	INVX1 INVX1_1971 ( .gnd(gnd), .vdd(vdd), .A(_11957_), .Y(_11958_) );
	NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_11958_), .B(_11954_), .Y(_11959_) );
	INVX1 INVX1_1972 ( .gnd(gnd), .vdd(vdd), .A(_11959_), .Y(_11960_) );
	NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_11958_), .B(_11954_), .Y(_11961_) );
	AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_11960_), .B(_11961_), .Y(_11962_) );
	XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_11950_), .B(_11962_), .Y(_11963_) );
	AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_11963_), .B(_13489_), .Y(_11964_) );
	NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_28_), .B(_13687__bF_buf7), .Y(_11965_) );
	OAI21X1 OAI21X1_4923 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_13687__bF_buf6), .C(_11965_), .Y(_11966_) );
	OAI21X1 OAI21X1_4924 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_13470__bF_buf0), .C(_11412__bF_buf2), .Y(_11967_) );
	AOI21X1 AOI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_11967_), .C(_13464__bF_buf0), .Y(_11968_) );
	OAI21X1 OAI21X1_4925 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_11967_), .C(_11968_), .Y(_11969_) );
	OAI21X1 OAI21X1_4926 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_13776__bF_buf3), .C(_11969_), .Y(_11970_) );
	AOI21X1 AOI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_11966_), .B(_13458__bF_buf7), .C(_11970_), .Y(_11971_) );
	NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf2), .B(_11971_), .Y(_11972_) );
	INVX1 INVX1_1973 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_28_), .Y(_11973_) );
	AOI21X1 AOI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_11973_), .B(_13397__bF_buf0), .C(_13398__bF_buf2), .Y(_11974_) );
	OAI21X1 OAI21X1_4927 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_11972_), .C(_11974_), .Y(_11975_) );
	NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_13695__bF_buf3), .Y(_11976_) );
	AOI21X1 AOI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_11976_), .B(_13694__bF_buf2), .C(_13391__bF_buf5), .Y(_11977_) );
	OAI21X1 OAI21X1_4928 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_28_), .B(_13392__bF_buf0), .C(_13412__bF_buf1), .Y(_11978_) );
	AOI21X1 AOI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_11975_), .B(_11977_), .C(_11978_), .Y(_11293__28_) );
	NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_11962_), .B(_11950_), .Y(_11979_) );
	OAI21X1 OAI21X1_4929 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_11958_), .C(_11979_), .Y(_11980_) );
	INVX1 INVX1_1974 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_29_), .Y(_11981_) );
	OAI21X1 OAI21X1_4930 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf6), .B(_13466__bF_buf6), .C(biu_biu_data_out_29_), .Y(_11982_) );
	OAI21X1 OAI21X1_4931 ( .gnd(gnd), .vdd(vdd), .A(_11981_), .B(_13463__bF_buf1), .C(_11982_), .Y(_11983_) );
	INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .Y(_11984_) );
	OAI21X1 OAI21X1_4932 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(biu_pc_29_), .C(_11402__bF_buf1), .Y(_11985_) );
	OAI21X1 OAI21X1_4933 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13478__bF_buf2), .C(_11985_), .Y(_11986_) );
	INVX1 INVX1_1975 ( .gnd(gnd), .vdd(vdd), .A(_11986_), .Y(_11987_) );
	NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_11987_), .B(_11984_), .Y(_11988_) );
	INVX1 INVX1_1976 ( .gnd(gnd), .vdd(vdd), .A(_11988_), .Y(_11989_) );
	NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_11987_), .B(_11984_), .Y(_11990_) );
	NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_11990_), .B(_11989_), .Y(_11991_) );
	INVX1 INVX1_1977 ( .gnd(gnd), .vdd(vdd), .A(_11991_), .Y(_11992_) );
	OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_11980_), .B(_11992_), .Y(_11993_) );
	NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_11980_), .Y(_11994_) );
	NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_11994_), .B(_11993_), .Y(_11995_) );
	NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf0), .B(_11995_), .Y(_11996_) );
	NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_29_), .B(_13687__bF_buf5), .Y(_11997_) );
	OAI21X1 OAI21X1_4934 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13687__bF_buf4), .C(_11997_), .Y(_11998_) );
	OAI21X1 OAI21X1_4935 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .B(_13470__bF_buf4), .C(_11412__bF_buf1), .Y(_11999_) );
	AOI21X1 AOI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_11984_), .B(_11999_), .C(_13464__bF_buf3), .Y(_12000_) );
	OAI21X1 OAI21X1_4936 ( .gnd(gnd), .vdd(vdd), .A(_11984_), .B(_11999_), .C(_12000_), .Y(_12001_) );
	OAI21X1 OAI21X1_4937 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13776__bF_buf2), .C(_12001_), .Y(_12002_) );
	AOI21X1 AOI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_11998_), .B(_13458__bF_buf5), .C(_12002_), .Y(_12003_) );
	NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf1), .B(_12003_), .Y(_12004_) );
	INVX1 INVX1_1978 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_29_), .Y(_12005_) );
	AOI21X1 AOI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_12005_), .B(_13397__bF_buf4), .C(_13398__bF_buf1), .Y(_12006_) );
	OAI21X1 OAI21X1_4938 ( .gnd(gnd), .vdd(vdd), .A(_12004_), .B(_11996_), .C(_12006_), .Y(_12007_) );
	NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13695__bF_buf2), .Y(_12008_) );
	AOI21X1 AOI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_12008_), .B(_13694__bF_buf1), .C(_13391__bF_buf4), .Y(_12009_) );
	OAI21X1 OAI21X1_4939 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_29_), .B(_13392__bF_buf7), .C(_13412__bF_buf0), .Y(_12010_) );
	AOI21X1 AOI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_12007_), .B(_12009_), .C(_12010_), .Y(_11293__29_) );
	NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_11962_), .B(_11992_), .Y(_12011_) );
	INVX1 INVX1_1979 ( .gnd(gnd), .vdd(vdd), .A(_12011_), .Y(_12012_) );
	OAI21X1 OAI21X1_4940 ( .gnd(gnd), .vdd(vdd), .A(_11984_), .B(_11987_), .C(_11960_), .Y(_12013_) );
	AOI22X1 AOI22X1_660 ( .gnd(gnd), .vdd(vdd), .A(_11990_), .B(_12013_), .C(_12012_), .D(_11950_), .Y(_12014_) );
	INVX1 INVX1_1980 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_30_), .Y(_12015_) );
	OAI21X1 OAI21X1_4941 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf4), .B(_13466__bF_buf5), .C(biu_biu_data_out_30_), .Y(_12016_) );
	OAI21X1 OAI21X1_4942 ( .gnd(gnd), .vdd(vdd), .A(_12015_), .B(_13463__bF_buf0), .C(_12016_), .Y(_12017_) );
	OAI21X1 OAI21X1_4943 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(biu_pc_30_), .C(_11402__bF_buf0), .Y(_12018_) );
	OAI21X1 OAI21X1_4944 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13478__bF_buf1), .C(_12018_), .Y(_12019_) );
	XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .B(_12019_), .Y(_12020_) );
	AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_12014_), .B(_12020_), .Y(_12021_) );
	NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_12020_), .B(_12014_), .Y(_12022_) );
	NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12021_), .Y(_12023_) );
	NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf3), .B(_12023_), .Y(_12024_) );
	NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_30_), .B(_13687__bF_buf3), .Y(_12025_) );
	OAI21X1 OAI21X1_4945 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13687__bF_buf2), .C(_12025_), .Y(_12026_) );
	INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .Y(_12027_) );
	OAI21X1 OAI21X1_4946 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_13470__bF_buf3), .C(_11412__bF_buf0), .Y(_12028_) );
	AOI21X1 AOI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_12028_), .C(_13464__bF_buf2), .Y(_12029_) );
	OAI21X1 OAI21X1_4947 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_12028_), .C(_12029_), .Y(_12030_) );
	OAI21X1 OAI21X1_4948 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13776__bF_buf1), .C(_12030_), .Y(_12031_) );
	AOI21X1 AOI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_12026_), .B(_13458__bF_buf3), .C(_12031_), .Y(_12032_) );
	NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_13454__bF_buf0), .B(_12032_), .Y(_12033_) );
	INVX1 INVX1_1981 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_30_), .Y(_12034_) );
	AOI21X1 AOI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_12034_), .B(_13397__bF_buf3), .C(_13398__bF_buf0), .Y(_12035_) );
	OAI21X1 OAI21X1_4949 ( .gnd(gnd), .vdd(vdd), .A(_12024_), .B(_12033_), .C(_12035_), .Y(_12036_) );
	NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13695__bF_buf1), .Y(_12037_) );
	AOI21X1 AOI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_12037_), .B(_13694__bF_buf0), .C(_13391__bF_buf3), .Y(_12038_) );
	OAI21X1 OAI21X1_4950 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_30_), .B(_13392__bF_buf6), .C(_13412__bF_buf4), .Y(_12039_) );
	AOI21X1 AOI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_12036_), .B(_12038_), .C(_12039_), .Y(_11293__30_) );
	NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_12019_), .B(_12017_), .Y(_12040_) );
	NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_13971_), .B(_13972_), .C(_13825_), .Y(_12041_) );
	AOI21X1 AOI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_11502_), .B(_11508_), .C(_11551_), .Y(_12042_) );
	NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(_11479_), .B(_12042_), .C(_11445_), .Y(_12043_) );
	NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_12043_), .B(_11433_), .Y(_12044_) );
	OAI21X1 OAI21X1_4951 ( .gnd(gnd), .vdd(vdd), .A(_13977_), .B(_12041_), .C(_12044_), .Y(_12045_) );
	AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_11823_), .B(_11786_), .Y(_12046_) );
	NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(_11693_), .B(_11691_), .C(_12046_), .Y(_12047_) );
	AOI21X1 AOI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_12045_), .B(_11576_), .C(_12047_), .Y(_12048_) );
	NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_11895_), .B(_11946_), .Y(_12049_) );
	OAI21X1 OAI21X1_4952 ( .gnd(gnd), .vdd(vdd), .A(_11830_), .B(_12048_), .C(_12049_), .Y(_12050_) );
	AOI21X1 AOI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_12050_), .B(_11949_), .C(_12011_), .Y(_12051_) );
	OAI21X1 OAI21X1_4953 ( .gnd(gnd), .vdd(vdd), .A(_11960_), .B(_11991_), .C(_11989_), .Y(_12052_) );
	OAI21X1 OAI21X1_4954 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .B(_12051_), .C(_12020_), .Y(_12053_) );
	INVX1 INVX1_1982 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_31_), .Y(_12054_) );
	OAI21X1 OAI21X1_4955 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf2), .B(_13466__bF_buf4), .C(biu_biu_data_out_31_), .Y(_12055_) );
	OAI21X1 OAI21X1_4956 ( .gnd(gnd), .vdd(vdd), .A(_12054_), .B(_13463__bF_buf4), .C(_12055_), .Y(_12056_) );
	OAI21X1 OAI21X1_4957 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(biu_pc_31_), .C(_11402__bF_buf3), .Y(_12057_) );
	OAI21X1 OAI21X1_4958 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_13478__bF_buf0), .C(_12057_), .Y(_12058_) );
	XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .B(_12058_), .Y(_12059_) );
	INVX1 INVX1_1983 ( .gnd(gnd), .vdd(vdd), .A(_12059_), .Y(_12060_) );
	NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(_12040_), .B(_12060_), .C(_12053_), .Y(_12061_) );
	INVX1 INVX1_1984 ( .gnd(gnd), .vdd(vdd), .A(_12020_), .Y(_12062_) );
	OAI21X1 OAI21X1_4959 ( .gnd(gnd), .vdd(vdd), .A(_12062_), .B(_12014_), .C(_12040_), .Y(_12063_) );
	NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_12059_), .B(_12063_), .Y(_12064_) );
	NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_12061_), .B(_12064_), .Y(_12065_) );
	NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_13675_), .B(_13687__bF_buf1), .Y(_12066_) );
	OAI21X1 OAI21X1_4960 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_13687__bF_buf0), .C(_12066_), .Y(_12067_) );
	INVX1 INVX1_1985 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .Y(_12068_) );
	OAI21X1 OAI21X1_4961 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_13470__bF_buf2), .C(_11412__bF_buf3), .Y(_12069_) );
	OAI21X1 OAI21X1_4962 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12068_), .C(amoxor_bF_buf2), .Y(_12070_) );
	AOI21X1 AOI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_12068_), .B(_12069_), .C(_12070_), .Y(_12071_) );
	AOI21X1 AOI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(amoswap), .C(_12071_), .Y(_12072_) );
	OAI21X1 OAI21X1_4963 ( .gnd(gnd), .vdd(vdd), .A(_13459__bF_buf4), .B(_12067_), .C(_12072_), .Y(_12073_) );
	NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_12073_), .Y(_12074_) );
	OAI21X1 OAI21X1_4964 ( .gnd(gnd), .vdd(vdd), .A(_13488__bF_buf2), .B(_12065_), .C(_12074_), .Y(_12075_) );
	INVX1 INVX1_1986 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_31_), .Y(_12076_) );
	AOI21X1 AOI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_12076_), .B(_13397__bF_buf2), .C(_13398__bF_buf6), .Y(_12077_) );
	NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_12077_), .B(_12075_), .Y(_12078_) );
	NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_13695__bF_buf0), .Y(_12079_) );
	AOI21X1 AOI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_12079_), .B(_13694__bF_buf4), .C(_13391__bF_buf2), .Y(_12080_) );
	OAI21X1 OAI21X1_4965 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_in_31_), .B(_13392__bF_buf5), .C(_13412__bF_buf3), .Y(_12081_) );
	AOI21X1 AOI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_12078_), .B(_12080_), .C(_12081_), .Y(_11293__31_) );
	INVX1 INVX1_1987 ( .gnd(gnd), .vdd(vdd), .A(data_rd_0_), .Y(_12082_) );
	OAI21X1 OAI21X1_4966 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_13391__bF_buf1), .C(_13441__bF_buf3), .Y(_12083_) );
	INVX1 INVX1_1988 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltiu), .Y(_12084_) );
	OAI21X1 OAI21X1_4967 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_slti), .C(csr_gpr_iu_ins_dec_sltup), .Y(_12085_) );
	NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .Y(_12086_) );
	INVX4 INVX4_57 ( .gnd(gnd), .vdd(vdd), .A(_12086__bF_buf3), .Y(_12087_) );
	OAI21X1 OAI21X1_4968 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13640_), .Y(_12088_) );
	OAI21X1 OAI21X1_4969 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf3), .B(_12087_), .C(_12088_), .Y(_12089_) );
	OAI21X1 OAI21X1_4970 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .B(_13926_), .C(_12089_), .Y(_12090_) );
	OAI21X1 OAI21X1_4971 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13885_), .Y(_12091_) );
	OAI21X1 OAI21X1_4972 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf1), .B(_12087_), .C(_12091_), .Y(_12092_) );
	NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_13890_), .Y(_12093_) );
	INVX1 INVX1_1989 ( .gnd(gnd), .vdd(vdd), .A(_12093_), .Y(_12094_) );
	NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .B(_13944_), .Y(_12095_) );
	AOI21X1 AOI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_13890_), .B(_12092_), .C(_12095_), .Y(_12096_) );
	NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(_12090_), .B(_12094_), .C(_12096_), .Y(_12097_) );
	OAI21X1 OAI21X1_4973 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13612_), .Y(_12098_) );
	OAI21X1 OAI21X1_4974 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf3), .B(_12087_), .C(_12098_), .Y(_12099_) );
	NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_12099_), .B(_13856_), .Y(_12100_) );
	AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_13856_), .B(_12099_), .Y(_12101_) );
	NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_12100_), .B(_12101_), .Y(_12102_) );
	OAI21X1 OAI21X1_4975 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13451_), .Y(_12103_) );
	OAI21X1 OAI21X1_4976 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_4_), .B(_12087_), .C(_12103_), .Y(_12104_) );
	NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_12104_), .B(_13812_), .Y(_12105_) );
	AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_13812_), .B(_12104_), .Y(_12106_) );
	OAI21X1 OAI21X1_4977 ( .gnd(gnd), .vdd(vdd), .A(_12105_), .B(_12106_), .C(_12102_), .Y(_12107_) );
	NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_12107_), .B(_12097_), .Y(_12108_) );
	OAI21X1 OAI21X1_4978 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13435_), .Y(_12109_) );
	OAI21X1 OAI21X1_4979 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .B(_12087_), .C(_12109_), .Y(_12110_) );
	NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_12110_), .B(_13736_), .Y(_12111_) );
	OAI21X1 OAI21X1_4980 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_2_), .B(_13476__bF_buf3), .C(_13759_), .Y(_12112_) );
	OAI21X1 OAI21X1_4981 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13622_), .Y(_12113_) );
	OAI21X1 OAI21X1_4982 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_3_), .B(_12087_), .C(_12113_), .Y(_12114_) );
	XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_13779_), .B(_12114_), .Y(_12115_) );
	INVX1 INVX1_1990 ( .gnd(gnd), .vdd(vdd), .A(_12110_), .Y(_12116_) );
	OAI21X1 OAI21X1_4983 ( .gnd(gnd), .vdd(vdd), .A(_12112_), .B(_12116_), .C(_12115_), .Y(_12117_) );
	OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_12117_), .B(_12111_), .Y(_12118_) );
	OAI21X1 OAI21X1_4984 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13403_), .Y(_12119_) );
	OAI21X1 OAI21X1_4985 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(_12087_), .C(_12119_), .Y(_12120_) );
	OAI21X1 OAI21X1_4986 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13630_), .Y(_12121_) );
	OAI21X1 OAI21X1_4987 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_1_), .B(_12087_), .C(_12121_), .Y(_12122_) );
	NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .B(_13721_), .Y(_12123_) );
	INVX1 INVX1_1991 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .Y(_12124_) );
	INVX1 INVX1_1992 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .Y(_12125_) );
	NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_12120_), .B(_13468_), .Y(_12126_) );
	OAI21X1 OAI21X1_4988 ( .gnd(gnd), .vdd(vdd), .A(_12125_), .B(_12124_), .C(_12126_), .Y(_12127_) );
	NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_12123_), .B(_12127_), .Y(_12128_) );
	OAI21X1 OAI21X1_4989 ( .gnd(gnd), .vdd(vdd), .A(_13468_), .B(_12120_), .C(_12128_), .Y(_12129_) );
	NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12118_), .Y(_12130_) );
	INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(_11523_), .Y(_12131_) );
	NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_11401_), .B(_12086__bF_buf2), .Y(_12132_) );
	OAI21X1 OAI21X1_4990 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12133_) );
	OAI21X1 OAI21X1_4991 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_12086__bF_buf0), .C(_12132__bF_buf2), .Y(_12134_) );
	NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_12134_), .B(_11572_), .Y(_12135_) );
	AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_11572_), .B(_12134_), .Y(_12136_) );
	NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_12135_), .B(_12136_), .Y(_12137_) );
	OAI21X1 OAI21X1_4992 ( .gnd(gnd), .vdd(vdd), .A(_12131_), .B(_12133_), .C(_12137_), .Y(_12138_) );
	AOI21X1 AOI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_12131_), .B(_12133_), .C(_12138_), .Y(_12139_) );
	OAI21X1 OAI21X1_4993 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_12086__bF_buf3), .C(_12132__bF_buf1), .Y(_12140_) );
	INVX1 INVX1_1993 ( .gnd(gnd), .vdd(vdd), .A(_12140_), .Y(_12141_) );
	OAI21X1 OAI21X1_4994 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_12086__bF_buf2), .C(_12132__bF_buf0), .Y(_12142_) );
	NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_12142_), .B(_11437_), .Y(_12143_) );
	AOI21X1 AOI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_11484_), .B(_12141_), .C(_12143_), .Y(_12144_) );
	NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .B(_11484_), .Y(_12145_) );
	AOI21X1 AOI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_11437_), .B(_12142_), .C(_12145_), .Y(_12146_) );
	NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(_12144_), .B(_12146_), .C(_12139_), .Y(_12147_) );
	OAI21X1 OAI21X1_4995 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13596_), .Y(_12148_) );
	OAI21X1 OAI21X1_4996 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf1), .B(_12087_), .C(_12148_), .Y(_12149_) );
	NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_12149_), .B(_11332_), .Y(_12150_) );
	AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_11332_), .B(_12149_), .Y(_12151_) );
	NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_12150_), .B(_12151_), .Y(_12152_) );
	OAI21X1 OAI21X1_4997 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_13599_), .Y(_12153_) );
	OAI21X1 OAI21X1_4998 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf0), .B(_12087_), .C(_12153_), .Y(_12154_) );
	NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .B(_13964_), .Y(_12155_) );
	OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(_12154_), .Y(_12156_) );
	AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_12156_), .B(_12155_), .Y(_12157_) );
	OAI21X1 OAI21X1_4999 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_sltup), .C(_11351_), .Y(_12158_) );
	OAI21X1 OAI21X1_5000 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf3), .B(_12087_), .C(_12158_), .Y(_12159_) );
	NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_12159_), .B(_11373_), .Y(_12160_) );
	OAI21X1 OAI21X1_5001 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13476__bF_buf2), .C(_11398_), .Y(_12161_) );
	OAI21X1 OAI21X1_5002 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12162_) );
	OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_12161_), .B(_12162_), .Y(_12163_) );
	NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_12162_), .B(_12161_), .Y(_12164_) );
	OAI21X1 OAI21X1_5003 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11355_), .C(_12159_), .Y(_12165_) );
	NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(_12165_), .B(_12163_), .C(_12164_), .Y(_12166_) );
	NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_12160_), .B(_12166_), .Y(_12167_) );
	NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(_12152_), .B(_12157_), .C(_12167_), .Y(_12168_) );
	NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_12168_), .B(_12147_), .Y(_12169_) );
	NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(_12108_), .B(_12130_), .C(_12169_), .Y(_12170_) );
	OAI21X1 OAI21X1_5004 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_12086__bF_buf0), .C(_12132__bF_buf2), .Y(_12171_) );
	OAI21X1 OAI21X1_5005 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_12086__bF_buf3), .C(_12132__bF_buf1), .Y(_12172_) );
	AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .B(_12172_), .Y(_12173_) );
	NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_12172_), .B(_12056_), .Y(_12174_) );
	NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_12174_), .B(_12173_), .Y(_12175_) );
	OAI21X1 OAI21X1_5006 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .B(_12171_), .C(_12175_), .Y(_12176_) );
	AOI21X1 AOI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .B(_12171_), .C(_12176_), .Y(_12177_) );
	OAI21X1 OAI21X1_5007 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .B(_12086__bF_buf2), .C(_12132__bF_buf0), .Y(_12178_) );
	XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_12178_), .Y(_12179_) );
	OAI21X1 OAI21X1_5008 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12180_) );
	XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .B(_12180_), .Y(_12181_) );
	NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_12179_), .B(_12181_), .C(_12177_), .Y(_12182_) );
	OAI21X1 OAI21X1_5009 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .B(_12086__bF_buf0), .C(_12132__bF_buf2), .Y(_12183_) );
	NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_12183_), .B(_11834_), .Y(_12184_) );
	OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(_12183_), .Y(_12185_) );
	OAI21X1 OAI21X1_5010 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_12086__bF_buf3), .C(_12132__bF_buf1), .Y(_12186_) );
	NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .B(_11860_), .Y(_12187_) );
	AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(_12186_), .Y(_12188_) );
	NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_12187_), .B(_12188_), .Y(_12189_) );
	NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_12184_), .B(_12185_), .C(_12189_), .Y(_12190_) );
	OAI21X1 OAI21X1_5011 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_27_), .B(_12086__bF_buf2), .C(_12132__bF_buf0), .Y(_12191_) );
	NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_12191_), .B(_11921_), .Y(_12192_) );
	OAI21X1 OAI21X1_5012 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12193_) );
	NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_12193_), .B(_11886_), .Y(_12194_) );
	NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_12192_), .B(_12194_), .Y(_12195_) );
	NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_12191_), .B(_11921_), .Y(_12196_) );
	NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_12193_), .B(_11886_), .Y(_12197_) );
	NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .B(_12197_), .C(_12195_), .Y(_12198_) );
	OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_12190_), .B(_12198_), .Y(_12199_) );
	NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_12199_), .B(_12182_), .Y(_12200_) );
	OAI21X1 OAI21X1_5013 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_12086__bF_buf0), .C(_12132__bF_buf2), .Y(_12201_) );
	OAI21X1 OAI21X1_5014 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_23_), .B(_12086__bF_buf3), .C(_12132__bF_buf1), .Y(_12202_) );
	NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_12202_), .B(_11799_), .Y(_12203_) );
	AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_12202_), .Y(_12204_) );
	NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_12203_), .B(_12204_), .Y(_12205_) );
	OAI21X1 OAI21X1_5015 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_12201_), .C(_12205_), .Y(_12206_) );
	AOI21X1 AOI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_12201_), .C(_12206_), .Y(_12207_) );
	OAI21X1 OAI21X1_5016 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_12086__bF_buf2), .C(_12132__bF_buf0), .Y(_12208_) );
	XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_12208_), .Y(_12209_) );
	OAI21X1 OAI21X1_5017 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12210_) );
	XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .B(_12210_), .Y(_12211_) );
	NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(_12209_), .B(_12211_), .C(_12207_), .Y(_12212_) );
	OAI21X1 OAI21X1_5018 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_12086__bF_buf0), .C(_12132__bF_buf2), .Y(_12213_) );
	NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_12213_), .B(_11606_), .Y(_12214_) );
	INVX1 INVX1_1994 ( .gnd(gnd), .vdd(vdd), .A(_12214_), .Y(_12215_) );
	OAI21X1 OAI21X1_5019 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(_12086__bF_buf3), .C(_12132__bF_buf1), .Y(_12216_) );
	OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_11580_), .B(_12216_), .Y(_12217_) );
	AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_12215_), .B(_12217_), .Y(_12218_) );
	AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_11606_), .B(_12213_), .Y(_12219_) );
	AOI21X1 AOI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_11580_), .B(_12216_), .C(_12219_), .Y(_12220_) );
	INVX1 INVX1_1995 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_19_), .Y(_12221_) );
	OAI21X1 OAI21X1_5020 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf1), .B(_13466__bF_buf3), .C(biu_biu_data_out_19_), .Y(_12222_) );
	OAI21X1 OAI21X1_5021 ( .gnd(gnd), .vdd(vdd), .A(_12221_), .B(_13463__bF_buf3), .C(_12222_), .Y(_12223_) );
	OAI21X1 OAI21X1_5022 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_12086__bF_buf2), .C(_12132__bF_buf0), .Y(_12224_) );
	OAI21X1 OAI21X1_5023 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_12086__bF_buf1), .C(_12132__bF_buf3), .Y(_12225_) );
	OAI22X1 OAI22X1_822 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .B(_12223_), .C(_11662_), .D(_12225_), .Y(_12226_) );
	INVX1 INVX1_1996 ( .gnd(gnd), .vdd(vdd), .A(_12225_), .Y(_12227_) );
	NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .B(_12223_), .Y(_12228_) );
	OAI21X1 OAI21X1_5024 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_12227_), .C(_12228_), .Y(_12229_) );
	NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_12229_), .B(_12226_), .Y(_12230_) );
	NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(_12220_), .B(_12218_), .C(_12230_), .Y(_12231_) );
	NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_12231_), .B(_12212_), .Y(_12232_) );
	NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12232_), .Y(_12233_) );
	INVX1 INVX1_1997 ( .gnd(gnd), .vdd(vdd), .A(_12123_), .Y(_12234_) );
	AOI21X1 AOI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_12234_), .B(_12127_), .C(_12118_), .Y(_12235_) );
	OAI21X1 OAI21X1_5025 ( .gnd(gnd), .vdd(vdd), .A(_13624_), .B(_13476__bF_buf1), .C(_13786_), .Y(_12236_) );
	NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_12111_), .B(_12115_), .Y(_12237_) );
	OAI21X1 OAI21X1_5026 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .B(_12114_), .C(_12237_), .Y(_12238_) );
	OAI21X1 OAI21X1_5027 ( .gnd(gnd), .vdd(vdd), .A(_12238_), .B(_12235_), .C(_12108_), .Y(_12239_) );
	NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_12104_), .B(_13863_), .Y(_12240_) );
	AOI21X1 AOI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_12102_), .B(_12240_), .C(_12100_), .Y(_12241_) );
	OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_12097_), .B(_12241_), .Y(_12242_) );
	AOI21X1 AOI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_12090_), .B(_12093_), .C(_12095_), .Y(_12243_) );
	NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(_12242_), .B(_12243_), .C(_12239_), .Y(_12244_) );
	NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_12145_), .B(_12144_), .Y(_12245_) );
	INVX1 INVX1_1998 ( .gnd(gnd), .vdd(vdd), .A(_12135_), .Y(_12246_) );
	OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_12131_), .B(_12133_), .Y(_12247_) );
	OAI21X1 OAI21X1_5028 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12247_), .C(_12246_), .Y(_12248_) );
	AOI21X1 AOI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_12139_), .B(_12245_), .C(_12248_), .Y(_12249_) );
	INVX1 INVX1_1999 ( .gnd(gnd), .vdd(vdd), .A(_12160_), .Y(_12250_) );
	OAI21X1 OAI21X1_5029 ( .gnd(gnd), .vdd(vdd), .A(_12161_), .B(_12162_), .C(_12250_), .Y(_12251_) );
	INVX1 INVX1_2000 ( .gnd(gnd), .vdd(vdd), .A(_12150_), .Y(_12252_) );
	OAI21X1 OAI21X1_5030 ( .gnd(gnd), .vdd(vdd), .A(_12156_), .B(_12151_), .C(_12252_), .Y(_12253_) );
	AOI22X1 AOI22X1_661 ( .gnd(gnd), .vdd(vdd), .A(_12167_), .B(_12253_), .C(_12164_), .D(_12251_), .Y(_12254_) );
	OAI21X1 OAI21X1_5031 ( .gnd(gnd), .vdd(vdd), .A(_12254_), .B(_12147_), .C(_12249_), .Y(_12255_) );
	AOI21X1 AOI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_12244_), .B(_12169_), .C(_12255_), .Y(_12256_) );
	NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_12180_), .B(_11953_), .Y(_12257_) );
	NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_12257_), .B(_12179_), .Y(_12258_) );
	OAI21X1 OAI21X1_5032 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_12178_), .C(_12258_), .Y(_12259_) );
	INVX1 INVX1_2001 ( .gnd(gnd), .vdd(vdd), .A(_12174_), .Y(_12260_) );
	OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .B(_12171_), .Y(_12261_) );
	OAI21X1 OAI21X1_5033 ( .gnd(gnd), .vdd(vdd), .A(_12261_), .B(_12173_), .C(_12260_), .Y(_12262_) );
	AOI21X1 AOI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_12177_), .B(_12259_), .C(_12262_), .Y(_12263_) );
	AOI21X1 AOI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .B(_12191_), .C(_12195_), .Y(_12264_) );
	NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_12188_), .B(_12185_), .Y(_12265_) );
	NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_12187_), .B(_12265_), .Y(_12266_) );
	NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_12198_), .B(_12266_), .Y(_12267_) );
	NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_12264_), .B(_12267_), .Y(_12268_) );
	OAI21X1 OAI21X1_5034 ( .gnd(gnd), .vdd(vdd), .A(_12182_), .B(_12268_), .C(_12263_), .Y(_12269_) );
	OAI21X1 OAI21X1_5035 ( .gnd(gnd), .vdd(vdd), .A(_12217_), .B(_12219_), .C(_12215_), .Y(_12270_) );
	AOI22X1 AOI22X1_662 ( .gnd(gnd), .vdd(vdd), .A(_12226_), .B(_12228_), .C(_12270_), .D(_12230_), .Y(_12271_) );
	NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_12210_), .B(_11698_), .Y(_12272_) );
	NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .B(_12209_), .Y(_12273_) );
	OAI21X1 OAI21X1_5036 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_12208_), .C(_12273_), .Y(_12274_) );
	INVX1 INVX1_2002 ( .gnd(gnd), .vdd(vdd), .A(_12203_), .Y(_12275_) );
	OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_12201_), .Y(_12276_) );
	OAI21X1 OAI21X1_5037 ( .gnd(gnd), .vdd(vdd), .A(_12276_), .B(_12204_), .C(_12275_), .Y(_12277_) );
	AOI21X1 AOI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_12207_), .B(_12274_), .C(_12277_), .Y(_12278_) );
	OAI21X1 OAI21X1_5038 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .B(_12212_), .C(_12278_), .Y(_12279_) );
	AOI21X1 AOI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12279_), .C(_12269_), .Y(_12280_) );
	OAI21X1 OAI21X1_5039 ( .gnd(gnd), .vdd(vdd), .A(_12233_), .B(_12256_), .C(_12280_), .Y(_12281_) );
	OAI21X1 OAI21X1_5040 ( .gnd(gnd), .vdd(vdd), .A(_12170_), .B(_12233_), .C(_12281_), .Y(_12282_) );
	NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_sltp), .B(csr_gpr_iu_ins_dec_slti), .Y(_12283_) );
	NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_12283_), .B(_12173_), .Y(_12284_) );
	AOI22X1 AOI22X1_663 ( .gnd(gnd), .vdd(vdd), .A(_12084_), .B(_12085_), .C(_12284_), .D(_12282_), .Y(_12285_) );
	OAI21X1 OAI21X1_5041 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(addp_bF_buf2), .C(_13487_), .Y(_12286_) );
	NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13468_), .Y(_12287_) );
	NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf3), .B(_12287_), .Y(_12288_) );
	NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_orp), .B(csr_gpr_iu_ins_dec_ori), .Y(_12289_) );
	INVX8 INVX8_101 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .Y(_12290_) );
	NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .Y(_12291_) );
	MUX2X1 MUX2X1_169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(csr_gpr_iu_rs2_0_), .S(_12291__bF_buf3), .Y(_12292_) );
	NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_12292_), .B(_13469_), .Y(_12293_) );
	INVX4 INVX4_58 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf2), .Y(_12294_) );
	NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(andp), .B(andi), .Y(_12295_) );
	NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .Y(_12296_) );
	INVX8 INVX8_102 ( .gnd(gnd), .vdd(vdd), .A(_12296_), .Y(_12297_) );
	OAI21X1 OAI21X1_5042 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .C(_13403_), .Y(_12298_) );
	OAI21X1 OAI21X1_5043 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(_12297__bF_buf4), .C(_12298_), .Y(_12299_) );
	OAI22X1 OAI22X1_823 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_12294_), .C(_12295_), .D(_12299_), .Y(_12300_) );
	NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_12300_), .B(_13468_), .Y(_12301_) );
	NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrsi), .B(csr_gpr_iu_csrrwi), .Y(_12302_) );
	NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrw), .B(csr_gpr_iu_csrrci), .Y(_12303_) );
	NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrc), .B(csr_gpr_iu_csrrs), .Y(_12304_) );
	NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12303_), .C(_12304_), .Y(_12305_) );
	NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_ins_dec_jal_bF_buf7), .Y(_12306_) );
	OAI21X1 OAI21X1_5044 ( .gnd(gnd), .vdd(vdd), .A(_13479_), .B(_12306_), .C(_13398__bF_buf5), .Y(_12307_) );
	AOI21X1 AOI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(csr_0_), .B(_12305__bF_buf4), .C(_12307_), .Y(_12308_) );
	NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(_13467_), .B(_12301_), .C(_12308_), .Y(_12309_) );
	AOI21X1 AOI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf4), .B(_12293_), .C(_12309_), .Y(_12310_) );
	NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(_12288_), .B(_12286_), .C(_12310_), .Y(_12311_) );
	OAI21X1 OAI21X1_5045 ( .gnd(gnd), .vdd(vdd), .A(_12311_), .B(_12285_), .C(_12083_), .Y(_12312_) );
	NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(data_rd_1_), .B(_13416__bF_buf2), .Y(_12313_) );
	OAI21X1 OAI21X1_5046 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_13416__bF_buf1), .C(_12313_), .Y(_12314_) );
	NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(_13414_), .B(_13391__bF_buf0), .C(_12314_), .Y(_12315_) );
	AOI21X1 AOI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_12312_), .B(_12315_), .C(rst_bF_buf10), .Y(_11292__0_) );
	INVX1 INVX1_2003 ( .gnd(gnd), .vdd(vdd), .A(data_rd_1_), .Y(_12316_) );
	INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(data_rd_2_), .Y(_12317_) );
	MUX2X1 MUX2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12316_), .S(_13416__bF_buf0), .Y(_12318_) );
	AOI21X1 AOI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_13415__bF_buf4), .C(_13392__bF_buf4), .Y(_12319_) );
	OAI21X1 OAI21X1_5047 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf3), .B(_12318_), .C(_12319_), .Y(_12320_) );
	NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_12316_), .B(_13398__bF_buf4), .Y(_12321_) );
	INVX1 INVX1_2004 ( .gnd(gnd), .vdd(vdd), .A(_12287_), .Y(_12322_) );
	NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(_13721_), .Y(_12323_) );
	INVX1 INVX1_2005 ( .gnd(gnd), .vdd(vdd), .A(_12323_), .Y(_12324_) );
	NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(_13721_), .Y(_12325_) );
	NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_12325_), .B(_12324_), .Y(_12326_) );
	AOI21X1 AOI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_12326_), .B(_12322_), .C(_12294_), .Y(_12327_) );
	OAI21X1 OAI21X1_5048 ( .gnd(gnd), .vdd(vdd), .A(_12322_), .B(_12326_), .C(_12327_), .Y(_12328_) );
	INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(_12295_), .Y(_12329_) );
	OAI21X1 OAI21X1_5049 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(_12296_), .C(_12329_), .Y(_12330_) );
	AOI21X1 AOI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_13708_), .B(_12296_), .C(_12330_), .Y(_12331_) );
	OAI21X1 OAI21X1_5050 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(addp_bF_buf1), .C(_13719_), .Y(_12332_) );
	INVX8 INVX8_103 ( .gnd(gnd), .vdd(vdd), .A(_12291__bF_buf2), .Y(_12333_) );
	OAI21X1 OAI21X1_5051 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(csr_gpr_iu_rs2_1_), .Y(_12334_) );
	OAI21X1 OAI21X1_5052 ( .gnd(gnd), .vdd(vdd), .A(_13708_), .B(_12333_), .C(_12334_), .Y(_12335_) );
	OAI21X1 OAI21X1_5053 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(_13721_), .C(_12290__bF_buf3), .Y(_12336_) );
	INVX8 INVX8_104 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .Y(_12337_) );
	AOI22X1 AOI22X1_664 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .B(_12337__bF_buf3), .C(csr_1_), .D(_12305__bF_buf3), .Y(_12338_) );
	AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_12338_), .B(_13714_), .Y(_12339_) );
	NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(_12336_), .B(_12339_), .C(_12332_), .Y(_12340_) );
	AOI21X1 AOI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .B(_12331_), .C(_12340_), .Y(_12341_) );
	AOI21X1 AOI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .B(_12328_), .C(_13695__bF_buf5), .Y(_12342_) );
	OAI21X1 OAI21X1_5054 ( .gnd(gnd), .vdd(vdd), .A(_12321_), .B(_12342_), .C(_13392__bF_buf3), .Y(_12343_) );
	AOI21X1 AOI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_12343_), .B(_12320_), .C(rst_bF_buf9), .Y(_11292__1_) );
	INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(data_rd_3_), .Y(_12344_) );
	MUX2X1 MUX2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_12344_), .B(_12317_), .S(_13416__bF_buf4), .Y(_12345_) );
	AOI21X1 AOI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_12316_), .B(_13415__bF_buf2), .C(_13392__bF_buf2), .Y(_12346_) );
	OAI21X1 OAI21X1_5055 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf1), .B(_12345_), .C(_12346_), .Y(_12347_) );
	NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(addp_bF_buf0), .Y(_12348_) );
	OAI21X1 OAI21X1_5056 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13435_), .Y(_12349_) );
	OAI21X1 OAI21X1_5057 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .B(_12333_), .C(_12349_), .Y(_12350_) );
	NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_12350_), .B(_12112_), .Y(_12351_) );
	AOI21X1 AOI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_12297__bF_buf3), .B(_13435_), .C(_12295_), .Y(_12352_) );
	OAI21X1 OAI21X1_5058 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .B(_12297__bF_buf2), .C(_12352_), .Y(_12353_) );
	AOI22X1 AOI22X1_665 ( .gnd(gnd), .vdd(vdd), .A(_13750_), .B(_12337__bF_buf2), .C(csr_2_), .D(_12305__bF_buf2), .Y(_12354_) );
	AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_12354_), .B(_13749_), .Y(_12355_) );
	OAI21X1 OAI21X1_5059 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .B(_12112_), .C(_12355_), .Y(_12356_) );
	AOI21X1 AOI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf2), .B(_12351_), .C(_12356_), .Y(_12357_) );
	OAI21X1 OAI21X1_5060 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_13763_), .C(_12357_), .Y(_12358_) );
	OAI21X1 OAI21X1_5061 ( .gnd(gnd), .vdd(vdd), .A(_12287_), .B(_12325_), .C(_12323_), .Y(_12359_) );
	INVX1 INVX1_2006 ( .gnd(gnd), .vdd(vdd), .A(_12359_), .Y(_12360_) );
	NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .B(_13736_), .Y(_12361_) );
	NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_12112_), .Y(_12362_) );
	NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_12361_), .B(_12362_), .Y(_12363_) );
	INVX1 INVX1_2007 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .Y(_12364_) );
	NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_12364_), .B(_12360_), .Y(_12365_) );
	OAI21X1 OAI21X1_5062 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12359_), .C(csr_gpr_iu_ins_dec_subp_bF_buf1), .Y(_12366_) );
	OAI21X1 OAI21X1_5063 ( .gnd(gnd), .vdd(vdd), .A(_12366_), .B(_12365_), .C(_13398__bF_buf3), .Y(_12367_) );
	OAI21X1 OAI21X1_5064 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_13391__bF_buf7), .C(_13441__bF_buf2), .Y(_12368_) );
	OAI21X1 OAI21X1_5065 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12367_), .C(_12368_), .Y(_12369_) );
	AOI21X1 AOI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .B(_12347_), .C(rst_bF_buf8), .Y(_11292__2_) );
	INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(data_rd_4_), .Y(_12370_) );
	MUX2X1 MUX2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_12344_), .S(_13416__bF_buf3), .Y(_12371_) );
	AOI21X1 AOI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_13415__bF_buf0), .C(_13392__bF_buf1), .Y(_12372_) );
	OAI21X1 OAI21X1_5066 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf6), .B(_12371_), .C(_12372_), .Y(_12373_) );
	NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_12344_), .B(_13398__bF_buf2), .Y(_12374_) );
	NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13736_), .Y(_12375_) );
	OAI21X1 OAI21X1_5067 ( .gnd(gnd), .vdd(vdd), .A(_12364_), .B(_12360_), .C(_12375_), .Y(_12376_) );
	NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .B(_12236_), .Y(_12377_) );
	NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_13779_), .Y(_12378_) );
	NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_12377_), .B(_12378_), .Y(_12379_) );
	AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_12376_), .B(_12379_), .Y(_12380_) );
	OAI21X1 OAI21X1_5068 ( .gnd(gnd), .vdd(vdd), .A(_12379_), .B(_12376_), .C(csr_gpr_iu_ins_dec_subp_bF_buf0), .Y(_12381_) );
	INVX1 INVX1_2008 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_3_), .Y(_12382_) );
	OAI21X1 OAI21X1_5069 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .B(_12296_), .C(_12329_), .Y(_12383_) );
	AOI21X1 AOI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_12382_), .B(_12296_), .C(_12383_), .Y(_12384_) );
	OAI21X1 OAI21X1_5070 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(addp_bF_buf4), .C(_13800_), .Y(_12385_) );
	OAI21X1 OAI21X1_5071 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(csr_gpr_iu_rs2_3_), .Y(_12386_) );
	OAI21X1 OAI21X1_5072 ( .gnd(gnd), .vdd(vdd), .A(_12382_), .B(_12333_), .C(_12386_), .Y(_12387_) );
	OAI21X1 OAI21X1_5073 ( .gnd(gnd), .vdd(vdd), .A(_12387_), .B(_12236_), .C(_12290__bF_buf1), .Y(_12388_) );
	OAI21X1 OAI21X1_5074 ( .gnd(gnd), .vdd(vdd), .A(_13750_), .B(_13787_), .C(_12337__bF_buf1), .Y(_12389_) );
	AOI21X1 AOI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_13750_), .B(_13787_), .C(_12389_), .Y(_12390_) );
	INVX1 INVX1_2009 ( .gnd(gnd), .vdd(vdd), .A(csr_3_), .Y(_12391_) );
	INVX1 INVX1_2010 ( .gnd(gnd), .vdd(vdd), .A(_12305__bF_buf1), .Y(_12392_) );
	OAI21X1 OAI21X1_5075 ( .gnd(gnd), .vdd(vdd), .A(_12391_), .B(_12392_), .C(_13785_), .Y(_12393_) );
	NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_12390_), .B(_12393_), .Y(_12394_) );
	NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12394_), .C(_12385_), .Y(_12395_) );
	AOI21X1 AOI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .B(_12384_), .C(_12395_), .Y(_12396_) );
	OAI21X1 OAI21X1_5076 ( .gnd(gnd), .vdd(vdd), .A(_12380_), .B(_12381_), .C(_12396_), .Y(_12397_) );
	AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_12397_), .B(_13398__bF_buf1), .Y(_12398_) );
	OAI21X1 OAI21X1_5077 ( .gnd(gnd), .vdd(vdd), .A(_12374_), .B(_12398_), .C(_13392__bF_buf0), .Y(_12399_) );
	AOI21X1 AOI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12373_), .C(rst_bF_buf7), .Y(_11292__3_) );
	INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(data_rd_5_), .Y(_12400_) );
	MUX2X1 MUX2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_12400_), .B(_12370_), .S(_13416__bF_buf2), .Y(_12401_) );
	AOI21X1 AOI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_12344_), .B(_13415__bF_buf5), .C(_13392__bF_buf7), .Y(_12402_) );
	OAI21X1 OAI21X1_5078 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf4), .B(_12401_), .C(_12402_), .Y(_12403_) );
	OAI21X1 OAI21X1_5079 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_13391__bF_buf6), .C(_13441__bF_buf1), .Y(_12404_) );
	INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .Y(_12405_) );
	AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_13845_), .B(_12405_), .Y(_12406_) );
	NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(_13451_), .B(_13836_), .C(_13811_), .Y(_12407_) );
	NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_4_), .B(_13826_), .C(_13827_), .Y(_12408_) );
	NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_12407_), .B(_12408_), .Y(_12409_) );
	NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_12236_), .Y(_12410_) );
	NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_12236_), .Y(_12411_) );
	OAI21X1 OAI21X1_5080 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12411_), .C(_12410_), .Y(_12412_) );
	AOI22X1 AOI22X1_666 ( .gnd(gnd), .vdd(vdd), .A(_12361_), .B(_12362_), .C(_12377_), .D(_12378_), .Y(_12413_) );
	AOI21X1 AOI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_12359_), .B(_12413_), .C(_12412_), .Y(_12414_) );
	AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_12414_), .B(_12409_), .Y(_12415_) );
	OAI21X1 OAI21X1_5081 ( .gnd(gnd), .vdd(vdd), .A(_12409_), .B(_12414_), .C(csr_gpr_iu_ins_dec_subp_bF_buf3), .Y(_12416_) );
	OAI21X1 OAI21X1_5082 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_4_), .B(_12296_), .C(_12329_), .Y(_12417_) );
	AOI21X1 AOI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_13813_), .B(_12296_), .C(_12417_), .Y(_12418_) );
	OAI21X1 OAI21X1_5083 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13451_), .Y(_12419_) );
	OAI21X1 OAI21X1_5084 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_4_), .B(_12333_), .C(_12419_), .Y(_12420_) );
	AOI21X1 AOI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_13827_), .B(_12420_), .C(_12289_), .Y(_12421_) );
	NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(csr_4_), .B(_12305__bF_buf0), .Y(_12422_) );
	OAI21X1 OAI21X1_5085 ( .gnd(gnd), .vdd(vdd), .A(_13750_), .B(_13787_), .C(_13828_), .Y(_12423_) );
	NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_2_), .B(biu_pc_3_), .C(biu_pc_4_), .Y(_12424_) );
	AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf0), .B(_12424_), .Y(_12425_) );
	AOI21X1 AOI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_12423_), .B(_12425_), .C(_13695__bF_buf4), .Y(_12426_) );
	NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(_13826_), .B(_12422_), .C(_12426_), .Y(_12427_) );
	OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_12427_), .B(_12421_), .Y(_12428_) );
	AOI21X1 AOI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_13863_), .B(_12418_), .C(_12428_), .Y(_12429_) );
	OAI21X1 OAI21X1_5086 ( .gnd(gnd), .vdd(vdd), .A(_12415_), .B(_12416_), .C(_12429_), .Y(_12430_) );
	OAI21X1 OAI21X1_5087 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .B(_12430_), .C(_12404_), .Y(_12431_) );
	AOI21X1 AOI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_12431_), .B(_12403_), .C(rst_bF_buf6), .Y(_11292__4_) );
	INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(data_rd_6_), .Y(_12432_) );
	MUX2X1 MUX2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_12432_), .B(_12400_), .S(_13416__bF_buf1), .Y(_12433_) );
	AOI21X1 AOI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_13415__bF_buf3), .C(_13392__bF_buf6), .Y(_12434_) );
	OAI21X1 OAI21X1_5088 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf2), .B(_12433_), .C(_12434_), .Y(_12435_) );
	OAI21X1 OAI21X1_5089 ( .gnd(gnd), .vdd(vdd), .A(_12400_), .B(_13391__bF_buf5), .C(_13441__bF_buf0), .Y(_12436_) );
	NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_13877_), .Y(_12437_) );
	NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(_13612_), .B(_13865_), .C(_13866_), .Y(_12438_) );
	NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_5_), .B(_13855_), .C(_13874_), .Y(_12439_) );
	NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_12438_), .B(_12439_), .Y(_12440_) );
	INVX1 INVX1_2011 ( .gnd(gnd), .vdd(vdd), .A(_12440_), .Y(_12441_) );
	OAI21X1 OAI21X1_5090 ( .gnd(gnd), .vdd(vdd), .A(_12409_), .B(_12414_), .C(_12407_), .Y(_12442_) );
	AOI21X1 AOI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_12442_), .B(_12441_), .C(_12294_), .Y(_12443_) );
	OAI21X1 OAI21X1_5091 ( .gnd(gnd), .vdd(vdd), .A(_12441_), .B(_12442_), .C(_12443_), .Y(_12444_) );
	OAI21X1 OAI21X1_5092 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13612_), .Y(_12445_) );
	OAI21X1 OAI21X1_5093 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf2), .B(_12333_), .C(_12445_), .Y(_12446_) );
	OAI21X1 OAI21X1_5094 ( .gnd(gnd), .vdd(vdd), .A(_13854_), .B(_13463__bF_buf2), .C(_12446_), .Y(_12447_) );
	OAI21X1 OAI21X1_5095 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_orp), .B(csr_gpr_iu_ins_dec_ori), .C(_12447_), .Y(_12448_) );
	AOI21X1 AOI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_12297__bF_buf1), .B(_13612_), .C(_12295_), .Y(_12449_) );
	OAI21X1 OAI21X1_5096 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf1), .B(_12297__bF_buf0), .C(_12449_), .Y(_12450_) );
	NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_12450_), .B(_13874_), .Y(_12451_) );
	AOI21X1 AOI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_12424_), .B(_13867_), .C(_12306_), .Y(_12452_) );
	OAI21X1 OAI21X1_5097 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_12424_), .C(_12452_), .Y(_12453_) );
	AOI21X1 AOI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(csr_5_), .B(_12305__bF_buf4), .C(_13695__bF_buf3), .Y(_12454_) );
	NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_12453_), .C(_12454_), .Y(_12455_) );
	NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_12451_), .B(_12455_), .Y(_12456_) );
	NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(_12448_), .B(_12456_), .C(_12444_), .Y(_12457_) );
	OAI21X1 OAI21X1_5098 ( .gnd(gnd), .vdd(vdd), .A(_12437_), .B(_12457_), .C(_12436_), .Y(_12458_) );
	AOI21X1 AOI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_12458_), .B(_12435_), .C(rst_bF_buf5), .Y(_11292__5_) );
	INVX2 INVX2_161 ( .gnd(gnd), .vdd(vdd), .A(data_rd_7_), .Y(_12459_) );
	MUX2X1 MUX2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_12459_), .B(_12432_), .S(_13416__bF_buf0), .Y(_12460_) );
	AOI21X1 AOI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_12400_), .B(_13415__bF_buf1), .C(_13392__bF_buf5), .Y(_12461_) );
	OAI21X1 OAI21X1_5099 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf0), .B(_12460_), .C(_12461_), .Y(_12462_) );
	NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_12441_), .B(_12442_), .Y(_12463_) );
	NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_12438_), .B(_12463_), .Y(_12464_) );
	INVX1 INVX1_2012 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .Y(_12465_) );
	NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_13890_), .Y(_12466_) );
	NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .B(_13920_), .Y(_12467_) );
	NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_12466_), .B(_12467_), .Y(_12468_) );
	OAI21X1 OAI21X1_5100 ( .gnd(gnd), .vdd(vdd), .A(_12468_), .B(_12465_), .C(csr_gpr_iu_ins_dec_subp_bF_buf2), .Y(_12469_) );
	AOI21X1 AOI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12468_), .C(_12469_), .Y(_12470_) );
	OAI21X1 OAI21X1_5101 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(addp_bF_buf3), .C(_13911_), .Y(_12471_) );
	OAI21X1 OAI21X1_5102 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_12424_), .C(_13897_), .Y(_12472_) );
	NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_5_), .B(biu_pc_6_), .Y(_12473_) );
	NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_12473_), .B(_12424_), .Y(_12474_) );
	INVX1 INVX1_2013 ( .gnd(gnd), .vdd(vdd), .A(_12474_), .Y(_12475_) );
	NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf3), .B(_12472_), .C(_12475_), .Y(_12476_) );
	OAI21X1 OAI21X1_5103 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13885_), .Y(_12477_) );
	OAI21X1 OAI21X1_5104 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf0), .B(_12333_), .C(_12477_), .Y(_12478_) );
	NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_12478_), .B(_13920_), .Y(_12479_) );
	AOI21X1 AOI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_12297__bF_buf4), .B(_13885_), .C(_12295_), .Y(_12480_) );
	OAI21X1 OAI21X1_5105 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf3), .B(_12297__bF_buf3), .C(_12480_), .Y(_12481_) );
	AOI22X1 AOI22X1_667 ( .gnd(gnd), .vdd(vdd), .A(csr_6_), .B(_12305__bF_buf3), .C(biu_biu_data_out_6_), .D(_13463__bF_buf1), .Y(_12482_) );
	OAI21X1 OAI21X1_5106 ( .gnd(gnd), .vdd(vdd), .A(_12481_), .B(_13920_), .C(_12482_), .Y(_12483_) );
	AOI21X1 AOI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf0), .B(_12479_), .C(_12483_), .Y(_12484_) );
	NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(_12476_), .B(_12484_), .C(_12471_), .Y(_12485_) );
	OAI21X1 OAI21X1_5107 ( .gnd(gnd), .vdd(vdd), .A(_12485_), .B(_12470_), .C(_13398__bF_buf0), .Y(_12486_) );
	OAI21X1 OAI21X1_5108 ( .gnd(gnd), .vdd(vdd), .A(_12432_), .B(_13398__bF_buf6), .C(_12486_), .Y(_12487_) );
	NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_13392__bF_buf4), .B(_12487_), .Y(_12488_) );
	AOI21X1 AOI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_12488_), .B(_12462_), .C(rst_bF_buf4), .Y(_11292__6_) );
	INVX2 INVX2_162 ( .gnd(gnd), .vdd(vdd), .A(data_rd_8_), .Y(_12489_) );
	MUX2X1 MUX2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_12489_), .B(_12459_), .S(_13416__bF_buf4), .Y(_12490_) );
	AOI21X1 AOI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_12432_), .B(_13415__bF_buf6), .C(_13392__bF_buf3), .Y(_12491_) );
	OAI21X1 OAI21X1_5109 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf5), .B(_12490_), .C(_12491_), .Y(_12492_) );
	OAI21X1 OAI21X1_5110 ( .gnd(gnd), .vdd(vdd), .A(_12468_), .B(_12465_), .C(_12466_), .Y(_12493_) );
	OAI21X1 OAI21X1_5111 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .B(_13926_), .C(csr_gpr_iu_rs2_7_), .Y(_12494_) );
	NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_13640_), .B(_13943_), .Y(_12495_) );
	NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_12494_), .B(_12495_), .Y(_12496_) );
	OAI21X1 OAI21X1_5112 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .B(_12493_), .C(csr_gpr_iu_ins_dec_subp_bF_buf1), .Y(_12497_) );
	AOI21X1 AOI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_12493_), .B(_12496_), .C(_12497_), .Y(_12498_) );
	OAI21X1 OAI21X1_5113 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(csr_gpr_iu_rs2_7_), .Y(_12499_) );
	OAI21X1 OAI21X1_5114 ( .gnd(gnd), .vdd(vdd), .A(_13945_), .B(_12333_), .C(_12499_), .Y(_12500_) );
	OAI21X1 OAI21X1_5115 ( .gnd(gnd), .vdd(vdd), .A(_12500_), .B(_13944_), .C(_12290__bF_buf4), .Y(_12501_) );
	NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf2), .B(_12296_), .Y(_12502_) );
	OAI21X1 OAI21X1_5116 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .C(csr_gpr_iu_rs2_7_), .Y(_12503_) );
	AOI21X1 AOI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_12502_), .B(_12503_), .C(_12295_), .Y(_12504_) );
	NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_13929_), .B(_12475_), .Y(_12505_) );
	INVX1 INVX1_2014 ( .gnd(gnd), .vdd(vdd), .A(_12505_), .Y(_12506_) );
	OAI21X1 OAI21X1_5117 ( .gnd(gnd), .vdd(vdd), .A(_12473_), .B(_12424_), .C(_13929_), .Y(_12507_) );
	NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf2), .B(_12507_), .C(_12506_), .Y(_12508_) );
	AOI21X1 AOI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(csr_7_), .B(_12305__bF_buf2), .C(_13695__bF_buf2), .Y(_12509_) );
	NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(_13925_), .B(_12508_), .C(_12509_), .Y(_12510_) );
	AOI21X1 AOI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_12504_), .C(_12510_), .Y(_12511_) );
	AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(_12511_), .B(_12501_), .Y(_12512_) );
	OAI21X1 OAI21X1_5118 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_13939_), .C(_12512_), .Y(_12513_) );
	OAI21X1 OAI21X1_5119 ( .gnd(gnd), .vdd(vdd), .A(_12459_), .B(_13391__bF_buf4), .C(_13441__bF_buf4), .Y(_12514_) );
	OAI21X1 OAI21X1_5120 ( .gnd(gnd), .vdd(vdd), .A(_12513_), .B(_12498_), .C(_12514_), .Y(_12515_) );
	AOI21X1 AOI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_12515_), .B(_12492_), .C(rst_bF_buf3), .Y(_11292__7_) );
	INVX2 INVX2_163 ( .gnd(gnd), .vdd(vdd), .A(data_rd_9_), .Y(_12516_) );
	MUX2X1 MUX2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_12516_), .B(_12489_), .S(_13416__bF_buf3), .Y(_12517_) );
	AOI21X1 AOI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_12459_), .B(_13415__bF_buf4), .C(_13392__bF_buf2), .Y(_12518_) );
	OAI21X1 OAI21X1_5121 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf3), .B(_12517_), .C(_12518_), .Y(_12519_) );
	XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(csr_gpr_iu_rs2_8_), .Y(_12520_) );
	OAI21X1 OAI21X1_5122 ( .gnd(gnd), .vdd(vdd), .A(_12407_), .B(_12440_), .C(_12438_), .Y(_12521_) );
	NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(_13943_), .Y(_12522_) );
	OAI21X1 OAI21X1_5123 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(_13943_), .C(_12466_), .Y(_12523_) );
	AOI21X1 AOI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_12494_), .B(_12495_), .C(_12468_), .Y(_12524_) );
	AOI22X1 AOI22X1_668 ( .gnd(gnd), .vdd(vdd), .A(_12522_), .B(_12523_), .C(_12521_), .D(_12524_), .Y(_12525_) );
	NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_12409_), .B(_12440_), .Y(_12526_) );
	NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_12526_), .B(_12524_), .Y(_12527_) );
	OAI21X1 OAI21X1_5124 ( .gnd(gnd), .vdd(vdd), .A(_12527_), .B(_12414_), .C(_12525_), .Y(_12528_) );
	NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_12520_), .B(_12528_), .Y(_12529_) );
	INVX1 INVX1_2015 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .Y(_12530_) );
	OAI21X1 OAI21X1_5125 ( .gnd(gnd), .vdd(vdd), .A(_12520_), .B(_12528_), .C(csr_gpr_iu_ins_dec_subp_bF_buf0), .Y(_12531_) );
	NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_12531_), .B(_12530_), .Y(_12532_) );
	OAI21X1 OAI21X1_5126 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(addp_bF_buf2), .C(_11302_), .Y(_12533_) );
	NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_13982_), .B(_12506_), .Y(_12534_) );
	INVX1 INVX1_2016 ( .gnd(gnd), .vdd(vdd), .A(_12534_), .Y(_12535_) );
	OAI21X1 OAI21X1_5127 ( .gnd(gnd), .vdd(vdd), .A(_13929_), .B(_12475_), .C(_13982_), .Y(_12536_) );
	NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf1), .B(_12536_), .C(_12535_), .Y(_12537_) );
	INVX1 INVX1_2017 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .Y(_12538_) );
	OAI21X1 OAI21X1_5128 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13599_), .Y(_12539_) );
	OAI21X1 OAI21X1_5129 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf3), .B(_12333_), .C(_12539_), .Y(_12540_) );
	NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_12540_), .B(_12538_), .Y(_12541_) );
	OAI21X1 OAI21X1_5130 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .C(csr_gpr_iu_rs2_8_), .Y(_12542_) );
	OAI21X1 OAI21X1_5131 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_12297__bF_buf2), .C(_12542_), .Y(_12543_) );
	NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(_12329_), .B(_12543_), .C(_13964_), .Y(_12544_) );
	NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(csr_8_), .B(_12305__bF_buf1), .Y(_12545_) );
	NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(_11299_), .B(_12545_), .C(_12544_), .Y(_12546_) );
	AOI21X1 AOI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf3), .B(_12541_), .C(_12546_), .Y(_12547_) );
	NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(_12537_), .B(_12547_), .C(_12533_), .Y(_12548_) );
	OAI21X1 OAI21X1_5132 ( .gnd(gnd), .vdd(vdd), .A(_12532_), .B(_12548_), .C(_13398__bF_buf5), .Y(_12549_) );
	OAI21X1 OAI21X1_5133 ( .gnd(gnd), .vdd(vdd), .A(_12489_), .B(_13398__bF_buf4), .C(_12549_), .Y(_12550_) );
	NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_13392__bF_buf1), .B(_12550_), .Y(_12551_) );
	AOI21X1 AOI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_12551_), .B(_12519_), .C(rst_bF_buf2), .Y(_11292__8_) );
	INVX2 INVX2_164 ( .gnd(gnd), .vdd(vdd), .A(data_rd_10_), .Y(_12552_) );
	MUX2X1 MUX2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_12552_), .B(_12516_), .S(_13416__bF_buf2), .Y(_12553_) );
	AOI21X1 AOI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_12489_), .B(_13415__bF_buf2), .C(_13392__bF_buf0), .Y(_12554_) );
	OAI21X1 OAI21X1_5134 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf1), .B(_12553_), .C(_12554_), .Y(_12555_) );
	OAI21X1 OAI21X1_5135 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_8_), .B(_12538_), .C(_12529_), .Y(_12556_) );
	OAI21X1 OAI21X1_5136 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .B(_11321_), .C(_13596_), .Y(_12557_) );
	INVX1 INVX1_2018 ( .gnd(gnd), .vdd(vdd), .A(_12557_), .Y(_12558_) );
	NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .B(_11332_), .Y(_12559_) );
	NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_12559_), .B(_12558_), .Y(_12560_) );
	AOI21X1 AOI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12560_), .C(_12294_), .Y(_12561_) );
	OAI21X1 OAI21X1_5137 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12560_), .C(_12561_), .Y(_12562_) );
	OAI21X1 OAI21X1_5138 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(addp_bF_buf1), .C(_11327_), .Y(_12563_) );
	NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .B(_11321_), .Y(_12564_) );
	OAI21X1 OAI21X1_5139 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_13596_), .Y(_12565_) );
	OAI21X1 OAI21X1_5140 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf0), .B(_12333_), .C(_12565_), .Y(_12566_) );
	NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_12566_), .B(_12564_), .Y(_12567_) );
	OAI21X1 OAI21X1_5141 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .C(csr_gpr_iu_rs2_9_), .Y(_12568_) );
	OAI21X1 OAI21X1_5142 ( .gnd(gnd), .vdd(vdd), .A(_11333_), .B(_12297__bF_buf1), .C(_12568_), .Y(_12569_) );
	OAI21X1 OAI21X1_5143 ( .gnd(gnd), .vdd(vdd), .A(andp), .B(andi), .C(_12569_), .Y(_12570_) );
	AOI21X1 AOI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(csr_9_), .B(_12305__bF_buf0), .C(_11321_), .Y(_12571_) );
	OAI21X1 OAI21X1_5144 ( .gnd(gnd), .vdd(vdd), .A(_12570_), .B(_12564_), .C(_12571_), .Y(_12572_) );
	AOI21X1 AOI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf2), .B(_12567_), .C(_12572_), .Y(_12573_) );
	NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(_12563_), .B(_12573_), .C(_12562_), .Y(_12574_) );
	NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_11315_), .B(_12534_), .Y(_12575_) );
	NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_9_), .B(_12535_), .Y(_12576_) );
	OAI21X1 OAI21X1_5145 ( .gnd(gnd), .vdd(vdd), .A(_12575_), .B(_12576_), .C(_12337__bF_buf0), .Y(_12577_) );
	NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf3), .B(_12577_), .Y(_12578_) );
	OAI21X1 OAI21X1_5146 ( .gnd(gnd), .vdd(vdd), .A(_12516_), .B(_13391__bF_buf3), .C(_13441__bF_buf3), .Y(_12579_) );
	OAI21X1 OAI21X1_5147 ( .gnd(gnd), .vdd(vdd), .A(_12578_), .B(_12574_), .C(_12579_), .Y(_12580_) );
	AOI21X1 AOI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_12580_), .B(_12555_), .C(rst_bF_buf1), .Y(_11292__9_) );
	INVX2 INVX2_165 ( .gnd(gnd), .vdd(vdd), .A(data_rd_11_), .Y(_12581_) );
	MUX2X1 MUX2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_12552_), .S(_13416__bF_buf1), .Y(_12582_) );
	AOI21X1 AOI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_12516_), .B(_13415__bF_buf0), .C(_13392__bF_buf7), .Y(_12583_) );
	OAI21X1 OAI21X1_5148 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf6), .B(_12582_), .C(_12583_), .Y(_12584_) );
	NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_12552_), .B(_13398__bF_buf2), .Y(_12585_) );
	OAI21X1 OAI21X1_5149 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11355_), .C(csr_gpr_iu_rs2_10_), .Y(_12586_) );
	NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_11351_), .B(_11372_), .Y(_12587_) );
	NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_12586_), .B(_12587_), .Y(_12588_) );
	INVX1 INVX1_2019 ( .gnd(gnd), .vdd(vdd), .A(_12588_), .Y(_12589_) );
	INVX1 INVX1_2020 ( .gnd(gnd), .vdd(vdd), .A(_12559_), .Y(_12590_) );
	AOI21X1 AOI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12590_), .C(_12558_), .Y(_12591_) );
	AOI21X1 AOI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_12591_), .B(_12589_), .C(_12294_), .Y(_12592_) );
	OAI21X1 OAI21X1_5150 ( .gnd(gnd), .vdd(vdd), .A(_12589_), .B(_12591_), .C(_12592_), .Y(_12593_) );
	NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_7_), .B(biu_pc_8_), .C(biu_pc_9_), .Y(_12594_) );
	INVX1 INVX1_2021 ( .gnd(gnd), .vdd(vdd), .A(_12594_), .Y(_12595_) );
	NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(_12595_), .C(_12474_), .Y(_12596_) );
	INVX1 INVX1_2022 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .Y(_12597_) );
	NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_12473_), .B(_12424_), .C(_12594_), .Y(_12598_) );
	OAI21X1 OAI21X1_5151 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(_12598_), .C(_12337__bF_buf3), .Y(_12599_) );
	NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_12597_), .B(_12599_), .Y(_12600_) );
	OAI21X1 OAI21X1_5152 ( .gnd(gnd), .vdd(vdd), .A(amoor), .B(csr_gpr_iu_ins_dec_orp), .C(_11351_), .Y(_12601_) );
	OAI21X1 OAI21X1_5153 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf2), .B(_12333_), .C(_12601_), .Y(_12602_) );
	NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_12602_), .B(_11372_), .Y(_12603_) );
	OAI21X1 OAI21X1_5154 ( .gnd(gnd), .vdd(vdd), .A(amoand), .B(andp), .C(csr_gpr_iu_rs2_10_), .Y(_12604_) );
	OAI21X1 OAI21X1_5155 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(_12297__bF_buf0), .C(_12604_), .Y(_12605_) );
	OAI21X1 OAI21X1_5156 ( .gnd(gnd), .vdd(vdd), .A(andp), .B(andi), .C(_12605_), .Y(_12606_) );
	AOI21X1 AOI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(csr_10_), .B(_12305__bF_buf4), .C(_11355_), .Y(_12607_) );
	OAI21X1 OAI21X1_5157 ( .gnd(gnd), .vdd(vdd), .A(_12606_), .B(_11372_), .C(_12607_), .Y(_12608_) );
	AOI21X1 AOI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf1), .B(_12603_), .C(_12608_), .Y(_12609_) );
	OAI21X1 OAI21X1_5158 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11368_), .C(_12609_), .Y(_12610_) );
	NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_12600_), .B(_12610_), .Y(_12611_) );
	AOI21X1 AOI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_12593_), .B(_12611_), .C(_13695__bF_buf1), .Y(_12612_) );
	OAI21X1 OAI21X1_5159 ( .gnd(gnd), .vdd(vdd), .A(_12585_), .B(_12612_), .C(_13392__bF_buf6), .Y(_12613_) );
	AOI21X1 AOI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12584_), .C(rst_bF_buf0), .Y(_11292__10_) );
	INVX2 INVX2_166 ( .gnd(gnd), .vdd(vdd), .A(data_rd_12_), .Y(_12614_) );
	MUX2X1 MUX2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_12614_), .B(_12581_), .S(_13416__bF_buf0), .Y(_12615_) );
	AOI21X1 AOI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_12552_), .B(_13415__bF_buf5), .C(_13392__bF_buf5), .Y(_12616_) );
	OAI21X1 OAI21X1_5160 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf4), .B(_12615_), .C(_12616_), .Y(_12617_) );
	OAI21X1 OAI21X1_5161 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11355_), .C(_11351_), .Y(_12618_) );
	OAI21X1 OAI21X1_5162 ( .gnd(gnd), .vdd(vdd), .A(_12589_), .B(_12591_), .C(_12618_), .Y(_12619_) );
	NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_12161_), .Y(_12620_) );
	NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .B(_11410_), .Y(_12621_) );
	NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12621_), .Y(_12622_) );
	AOI21X1 AOI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .B(_12622_), .C(_12294_), .Y(_12623_) );
	OAI21X1 OAI21X1_5163 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .B(_12622_), .C(_12623_), .Y(_12624_) );
	OAI21X1 OAI21X1_5164 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf5), .B(addp_bF_buf0), .C(_11406_), .Y(_12625_) );
	NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(_12333_), .Y(_12626_) );
	INVX1 INVX1_2023 ( .gnd(gnd), .vdd(vdd), .A(_12626_), .Y(_12627_) );
	OAI21X1 OAI21X1_5165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_12291__bF_buf1), .C(_12627_), .Y(_12628_) );
	NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .B(_11410_), .Y(_12629_) );
	OAI21X1 OAI21X1_5166 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(_12297__bF_buf4), .C(_12329_), .Y(_12630_) );
	INVX2 INVX2_167 ( .gnd(gnd), .vdd(vdd), .A(_12630_), .Y(_12631_) );
	OAI21X1 OAI21X1_5167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_12296_), .C(_12631_), .Y(_12632_) );
	AOI22X1 AOI22X1_669 ( .gnd(gnd), .vdd(vdd), .A(csr_11_), .B(_12305__bF_buf3), .C(biu_biu_data_out_11_), .D(_13463__bF_buf0), .Y(_12633_) );
	OAI21X1 OAI21X1_5168 ( .gnd(gnd), .vdd(vdd), .A(_12632_), .B(_11410_), .C(_12633_), .Y(_12634_) );
	AOI21X1 AOI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf0), .B(_12629_), .C(_12634_), .Y(_12635_) );
	NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(_12625_), .B(_12635_), .C(_12624_), .Y(_12636_) );
	NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_10_), .B(biu_pc_11_), .C(_12598_), .Y(_12637_) );
	INVX1 INVX1_2024 ( .gnd(gnd), .vdd(vdd), .A(_12637_), .Y(_12638_) );
	OAI21X1 OAI21X1_5169 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_11_), .B(_12597_), .C(_12337__bF_buf2), .Y(_12639_) );
	OAI21X1 OAI21X1_5170 ( .gnd(gnd), .vdd(vdd), .A(_12638_), .B(_12639_), .C(_13398__bF_buf1), .Y(_12640_) );
	OAI21X1 OAI21X1_5171 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_13391__bF_buf2), .C(_13441__bF_buf2), .Y(_12641_) );
	OAI21X1 OAI21X1_5172 ( .gnd(gnd), .vdd(vdd), .A(_12640_), .B(_12636_), .C(_12641_), .Y(_12642_) );
	AOI21X1 AOI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_12642_), .B(_12617_), .C(rst_bF_buf70), .Y(_11292__11_) );
	INVX2 INVX2_168 ( .gnd(gnd), .vdd(vdd), .A(data_rd_13_), .Y(_12643_) );
	MUX2X1 MUX2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_12643_), .B(_12614_), .S(_13416__bF_buf4), .Y(_12644_) );
	AOI21X1 AOI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_13415__bF_buf3), .C(_13392__bF_buf4), .Y(_12645_) );
	OAI21X1 OAI21X1_5173 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf2), .B(_12644_), .C(_12645_), .Y(_12646_) );
	OAI21X1 OAI21X1_5174 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_12291__bF_buf0), .C(_12627_), .Y(_12647_) );
	NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .B(_11454_), .Y(_12648_) );
	OAI21X1 OAI21X1_5175 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_12296_), .C(_12631_), .Y(_12649_) );
	INVX1 INVX1_2025 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .Y(_12650_) );
	NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_11399_), .B(_12650_), .C(_12596_), .Y(_12651_) );
	OAI21X1 OAI21X1_5176 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .B(_12638_), .C(_12337__bF_buf1), .Y(_12652_) );
	NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_12651_), .B(_12652_), .Y(_12653_) );
	AOI22X1 AOI22X1_670 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_12_), .C(csr_12_), .D(_12305__bF_buf2), .Y(_12654_) );
	OAI21X1 OAI21X1_5177 ( .gnd(gnd), .vdd(vdd), .A(_13580_), .B(_13476__bF_buf0), .C(_12654_), .Y(_12655_) );
	NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_12655_), .B(_12653_), .Y(_12656_) );
	OAI21X1 OAI21X1_5178 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_12649_), .C(_12656_), .Y(_12657_) );
	AOI21X1 AOI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf4), .B(_12648_), .C(_12657_), .Y(_12658_) );
	OAI21X1 OAI21X1_5179 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11450_), .C(_12658_), .Y(_12659_) );
	NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_13599_), .B(_13964_), .Y(_12660_) );
	OAI21X1 OAI21X1_5180 ( .gnd(gnd), .vdd(vdd), .A(_12660_), .B(_12559_), .C(_12557_), .Y(_12661_) );
	NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_11410_), .Y(_12662_) );
	AOI22X1 AOI22X1_671 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12621_), .C(_12586_), .D(_12587_), .Y(_12663_) );
	OAI21X1 OAI21X1_5181 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_11410_), .C(_12618_), .Y(_12664_) );
	AOI22X1 AOI22X1_672 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(_12664_), .C(_12661_), .D(_12663_), .Y(_12665_) );
	NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(_12520_), .B(_12560_), .C(_12663_), .Y(_12666_) );
	INVX1 INVX1_2026 ( .gnd(gnd), .vdd(vdd), .A(_12666_), .Y(_12667_) );
	NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_12667_), .B(_12528_), .Y(_12668_) );
	NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_12665_), .B(_12668_), .Y(_12669_) );
	NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_11437_), .Y(_12670_) );
	INVX1 INVX1_2027 ( .gnd(gnd), .vdd(vdd), .A(_12670_), .Y(_12671_) );
	NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_11437_), .Y(_12672_) );
	NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_12672_), .B(_12671_), .Y(_12673_) );
	AOI21X1 AOI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_12669_), .B(_12673_), .C(_12294_), .Y(_12674_) );
	OAI21X1 OAI21X1_5182 ( .gnd(gnd), .vdd(vdd), .A(_12669_), .B(_12673_), .C(_12674_), .Y(_12675_) );
	NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf0), .B(_12675_), .Y(_12676_) );
	OAI21X1 OAI21X1_5183 ( .gnd(gnd), .vdd(vdd), .A(_12614_), .B(_13391__bF_buf1), .C(_13441__bF_buf1), .Y(_12677_) );
	OAI21X1 OAI21X1_5184 ( .gnd(gnd), .vdd(vdd), .A(_12659_), .B(_12676_), .C(_12677_), .Y(_12678_) );
	AOI21X1 AOI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_12678_), .B(_12646_), .C(rst_bF_buf69), .Y(_11292__12_) );
	INVX2 INVX2_169 ( .gnd(gnd), .vdd(vdd), .A(data_rd_14_), .Y(_12679_) );
	MUX2X1 MUX2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_12643_), .S(_13416__bF_buf3), .Y(_12680_) );
	AOI21X1 AOI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_12614_), .B(_13415__bF_buf1), .C(_13392__bF_buf3), .Y(_12681_) );
	OAI21X1 OAI21X1_5185 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf0), .B(_12680_), .C(_12681_), .Y(_12682_) );
	OAI21X1 OAI21X1_5186 ( .gnd(gnd), .vdd(vdd), .A(_12643_), .B(_13391__bF_buf0), .C(_13441__bF_buf0), .Y(_12683_) );
	NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11480_), .Y(_12684_) );
	AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_12668_), .B(_12665_), .Y(_12685_) );
	OAI21X1 OAI21X1_5187 ( .gnd(gnd), .vdd(vdd), .A(_12672_), .B(_12685_), .C(_12670_), .Y(_12686_) );
	OAI21X1 OAI21X1_5188 ( .gnd(gnd), .vdd(vdd), .A(_11469_), .B(_13463__bF_buf4), .C(_11476_), .Y(_12687_) );
	NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_12687_), .Y(_12688_) );
	NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_11484_), .Y(_12689_) );
	AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_12688_), .B(_12689_), .Y(_12690_) );
	AOI21X1 AOI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_12686_), .B(_12690_), .C(_12294_), .Y(_12691_) );
	OAI21X1 OAI21X1_5189 ( .gnd(gnd), .vdd(vdd), .A(_12686_), .B(_12690_), .C(_12691_), .Y(_12692_) );
	NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_12650_), .B(_11471_), .C(_12637_), .Y(_12693_) );
	NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12693_), .Y(_12694_) );
	OAI21X1 OAI21X1_5190 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(_12651_), .C(_12694_), .Y(_12695_) );
	AOI21X1 AOI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_12297__bF_buf3), .C(_12630_), .Y(_12696_) );
	OAI21X1 OAI21X1_5191 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf3), .B(_12696_), .C(_12687_), .Y(_12697_) );
	NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .B(_12626_), .Y(_12698_) );
	OAI21X1 OAI21X1_5192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_12291__bF_buf3), .C(_12698_), .Y(_12699_) );
	NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(csr_13_), .B(_12305__bF_buf1), .Y(_12700_) );
	AOI21X1 AOI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_13_), .C(_13695__bF_buf0), .Y(_12701_) );
	NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(_12699_), .B(_12700_), .C(_12701_), .Y(_12702_) );
	AOI21X1 AOI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(biu_biu_data_out_13_), .B(_13463__bF_buf3), .C(_12702_), .Y(_12703_) );
	AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_12703_), .B(_12697_), .Y(_12704_) );
	NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(_12695_), .B(_12704_), .C(_12692_), .Y(_12705_) );
	OAI21X1 OAI21X1_5193 ( .gnd(gnd), .vdd(vdd), .A(_12684_), .B(_12705_), .C(_12683_), .Y(_12706_) );
	AOI21X1 AOI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_12706_), .B(_12682_), .C(rst_bF_buf68), .Y(_11292__13_) );
	INVX2 INVX2_170 ( .gnd(gnd), .vdd(vdd), .A(data_rd_15_), .Y(_12707_) );
	MUX2X1 MUX2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_12707_), .B(_12679_), .S(_13416__bF_buf2), .Y(_12708_) );
	AOI21X1 AOI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_12643_), .B(_13415__bF_buf6), .C(_13392__bF_buf2), .Y(_12709_) );
	OAI21X1 OAI21X1_5194 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf5), .B(_12708_), .C(_12709_), .Y(_12710_) );
	AOI21X1 AOI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_11519_), .B(_11516_), .C(_12348_), .Y(_12711_) );
	NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_11503_), .C(_11505_), .Y(_12712_) );
	NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_11523_), .Y(_12713_) );
	NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_12712_), .B(_12713_), .Y(_12714_) );
	INVX1 INVX1_2028 ( .gnd(gnd), .vdd(vdd), .A(_12689_), .Y(_12715_) );
	OAI21X1 OAI21X1_5195 ( .gnd(gnd), .vdd(vdd), .A(_12670_), .B(_12715_), .C(_12688_), .Y(_12716_) );
	INVX1 INVX1_2029 ( .gnd(gnd), .vdd(vdd), .A(_12716_), .Y(_12717_) );
	NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(_12673_), .B(_12690_), .C(_12669_), .Y(_12718_) );
	AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_12718_), .B(_12717_), .Y(_12719_) );
	NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_12714_), .B(_12719_), .Y(_12720_) );
	NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_12714_), .B(_12719_), .Y(_12721_) );
	NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf3), .B(_12721_), .Y(_12722_) );
	INVX1 INVX1_2030 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .Y(_12723_) );
	INVX1 INVX1_2031 ( .gnd(gnd), .vdd(vdd), .A(_12693_), .Y(_12724_) );
	NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(biu_pc_14_), .C(_12651_), .Y(_12725_) );
	OAI21X1 OAI21X1_5196 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_ins_dec_jal_bF_buf6), .C(_12725_), .Y(_12726_) );
	AOI21X1 AOI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_12723_), .B(_12724_), .C(_12726_), .Y(_12727_) );
	AOI21X1 AOI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_12297__bF_buf2), .C(_12630_), .Y(_12728_) );
	OAI21X1 OAI21X1_5197 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf2), .B(_12728_), .C(_12131_), .Y(_12729_) );
	OAI21X1 OAI21X1_5198 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_14_), .B(_12291__bF_buf2), .C(_12698_), .Y(_12730_) );
	NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(csr_14_), .B(_12305__bF_buf0), .Y(_12731_) );
	AOI21X1 AOI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_14_), .C(_13695__bF_buf5), .Y(_12732_) );
	NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(_12730_), .B(_12731_), .C(_12732_), .Y(_12733_) );
	INVX1 INVX1_2032 ( .gnd(gnd), .vdd(vdd), .A(_12733_), .Y(_12734_) );
	NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_12729_), .C(_12734_), .Y(_12735_) );
	NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_12727_), .B(_12735_), .Y(_12736_) );
	OAI21X1 OAI21X1_5199 ( .gnd(gnd), .vdd(vdd), .A(_12720_), .B(_12722_), .C(_12736_), .Y(_12737_) );
	OAI21X1 OAI21X1_5200 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_13391__bF_buf7), .C(_13441__bF_buf4), .Y(_12738_) );
	OAI21X1 OAI21X1_5201 ( .gnd(gnd), .vdd(vdd), .A(_12711_), .B(_12737_), .C(_12738_), .Y(_12739_) );
	AOI21X1 AOI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_12739_), .B(_12710_), .C(rst_bF_buf67), .Y(_11292__14_) );
	INVX2 INVX2_171 ( .gnd(gnd), .vdd(vdd), .A(data_rd_16_), .Y(_12740_) );
	MUX2X1 MUX2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_12740_), .B(_12707_), .S(_13416__bF_buf1), .Y(_12741_) );
	AOI21X1 AOI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_13415__bF_buf4), .C(_13392__bF_buf1), .Y(_12742_) );
	OAI21X1 OAI21X1_5202 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf3), .B(_12741_), .C(_12742_), .Y(_12743_) );
	OAI21X1 OAI21X1_5203 ( .gnd(gnd), .vdd(vdd), .A(_12707_), .B(_13391__bF_buf6), .C(_13441__bF_buf3), .Y(_12744_) );
	AOI21X1 AOI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_11550_), .B(_11552_), .C(_12348_), .Y(_12745_) );
	AOI21X1 AOI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_12131_), .C(_12720_), .Y(_12746_) );
	NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_11572_), .Y(_12747_) );
	NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_11556_), .Y(_12748_) );
	NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_12747_), .B(_12748_), .Y(_12749_) );
	AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_12746_), .B(_12749_), .Y(_12750_) );
	OAI21X1 OAI21X1_5204 ( .gnd(gnd), .vdd(vdd), .A(_12749_), .B(_12746_), .C(csr_gpr_iu_ins_dec_subp_bF_buf2), .Y(_12751_) );
	INVX1 INVX1_2033 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .Y(_12752_) );
	OAI21X1 OAI21X1_5205 ( .gnd(gnd), .vdd(vdd), .A(_12723_), .B(_12724_), .C(_12752_), .Y(_12753_) );
	NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(biu_pc_15_), .C(_12693_), .Y(_12754_) );
	AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_12754_), .B(_12337__bF_buf0), .Y(_12755_) );
	NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_11401_), .B(_12333_), .Y(_12756_) );
	INVX4 INVX4_59 ( .gnd(gnd), .vdd(vdd), .A(_12756_), .Y(_12757_) );
	OAI21X1 OAI21X1_5206 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_12291__bF_buf1), .C(_12757_), .Y(_12758_) );
	OAI21X1 OAI21X1_5207 ( .gnd(gnd), .vdd(vdd), .A(_12758_), .B(_11572_), .C(_12290__bF_buf1), .Y(_12759_) );
	AOI21X1 AOI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_12297__bF_buf1), .C(_12630_), .Y(_12760_) );
	NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(csr_15_), .B(_12305__bF_buf4), .Y(_12761_) );
	AOI21X1 AOI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_15_bF_buf4), .C(_13695__bF_buf4), .Y(_12762_) );
	NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(_11545_), .B(_12761_), .C(_12762_), .Y(_12763_) );
	AOI21X1 AOI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_11572_), .B(_12760_), .C(_12763_), .Y(_12764_) );
	NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_12759_), .B(_12764_), .Y(_12765_) );
	AOI21X1 AOI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_12755_), .B(_12753_), .C(_12765_), .Y(_12766_) );
	OAI21X1 OAI21X1_5208 ( .gnd(gnd), .vdd(vdd), .A(_12750_), .B(_12751_), .C(_12766_), .Y(_12767_) );
	OAI21X1 OAI21X1_5209 ( .gnd(gnd), .vdd(vdd), .A(_12745_), .B(_12767_), .C(_12744_), .Y(_12768_) );
	AOI21X1 AOI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_12768_), .B(_12743_), .C(rst_bF_buf66), .Y(_11292__15_) );
	INVX2 INVX2_172 ( .gnd(gnd), .vdd(vdd), .A(data_rd_17_), .Y(_12769_) );
	MUX2X1 MUX2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_12769_), .B(_12740_), .S(_13416__bF_buf0), .Y(_12770_) );
	AOI21X1 AOI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_12707_), .B(_13415__bF_buf2), .C(_13392__bF_buf0), .Y(_12771_) );
	OAI21X1 OAI21X1_5210 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf1), .B(_12770_), .C(_12771_), .Y(_12772_) );
	NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_12714_), .B(_12749_), .Y(_12773_) );
	NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(_12690_), .B(_12673_), .C(_12773_), .Y(_12774_) );
	NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_12666_), .B(_12774_), .Y(_12775_) );
	OAI21X1 OAI21X1_5211 ( .gnd(gnd), .vdd(vdd), .A(_12712_), .B(_12749_), .C(_12747_), .Y(_12776_) );
	AOI21X1 AOI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_12716_), .B(_12773_), .C(_12776_), .Y(_12777_) );
	OAI21X1 OAI21X1_5212 ( .gnd(gnd), .vdd(vdd), .A(_12665_), .B(_12774_), .C(_12777_), .Y(_12778_) );
	AOI21X1 AOI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_12775_), .B(_12528_), .C(_12778_), .Y(_12779_) );
	NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(_11589_), .Y(_12780_) );
	NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_11580_), .Y(_12781_) );
	OAI21X1 OAI21X1_5213 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_12781_), .C(_12779_), .Y(_12782_) );
	OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_12781_), .Y(_12783_) );
	OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_12779_), .B(_12783_), .Y(_12784_) );
	NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf1), .B(_12782_), .C(_12784_), .Y(_12785_) );
	OAI21X1 OAI21X1_5214 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf4), .B(addp_bF_buf4), .C(_11584_), .Y(_12786_) );
	AOI21X1 AOI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_12297__bF_buf0), .C(_12630_), .Y(_12787_) );
	AOI21X1 AOI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_12333_), .C(_12626_), .Y(_12788_) );
	OAI21X1 OAI21X1_5215 ( .gnd(gnd), .vdd(vdd), .A(_12788_), .B(_11580_), .C(_12290__bF_buf0), .Y(_12789_) );
	AOI22X1 AOI22X1_673 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_16_), .C(csr_16_), .D(_12305__bF_buf3), .Y(_12790_) );
	NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(_11579_), .B(_12790_), .C(_12789_), .Y(_12791_) );
	AOI21X1 AOI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_11580_), .B(_12787_), .C(_12791_), .Y(_12792_) );
	NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(_12792_), .B(_12785_), .C(_12786_), .Y(_12793_) );
	INVX2 INVX2_173 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .Y(_12794_) );
	AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_12754_), .B(_12794_), .Y(_12795_) );
	OAI21X1 OAI21X1_5216 ( .gnd(gnd), .vdd(vdd), .A(_12794_), .B(_12754_), .C(_12337__bF_buf3), .Y(_12796_) );
	OAI21X1 OAI21X1_5217 ( .gnd(gnd), .vdd(vdd), .A(_12796_), .B(_12795_), .C(_13398__bF_buf6), .Y(_12797_) );
	OAI21X1 OAI21X1_5218 ( .gnd(gnd), .vdd(vdd), .A(_12740_), .B(_13391__bF_buf5), .C(_13441__bF_buf2), .Y(_12798_) );
	OAI21X1 OAI21X1_5219 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .B(_12793_), .C(_12798_), .Y(_12799_) );
	AOI21X1 AOI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_12799_), .B(_12772_), .C(rst_bF_buf65), .Y(_11292__16_) );
	INVX2 INVX2_174 ( .gnd(gnd), .vdd(vdd), .A(data_rd_18_), .Y(_12800_) );
	MUX2X1 MUX2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_12769_), .S(_13416__bF_buf4), .Y(_12801_) );
	AOI21X1 AOI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_12740_), .B(_13415__bF_buf0), .C(_13392__bF_buf7), .Y(_12802_) );
	OAI21X1 OAI21X1_5220 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf6), .B(_12801_), .C(_12802_), .Y(_12803_) );
	OAI21X1 OAI21X1_5221 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf3), .B(addp_bF_buf3), .C(_11616_), .Y(_12804_) );
	NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12794_), .C(_12725_), .Y(_12805_) );
	INVX1 INVX1_2034 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .Y(_12806_) );
	NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_12794_), .B(_12806_), .C(_12754_), .Y(_12807_) );
	NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12807_), .Y(_12808_) );
	OAI21X1 OAI21X1_5222 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(_12805_), .C(_12808_), .Y(_12809_) );
	AOI21X1 AOI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_12297__bF_buf4), .C(_12630_), .Y(_12810_) );
	AOI21X1 AOI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_12333_), .C(_12626_), .Y(_12811_) );
	OAI21X1 OAI21X1_5223 ( .gnd(gnd), .vdd(vdd), .A(_12811_), .B(_11606_), .C(_12290__bF_buf4), .Y(_12812_) );
	AOI22X1 AOI22X1_674 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_17_), .C(csr_17_), .D(_12305__bF_buf2), .Y(_12813_) );
	NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(_11605_), .B(_12813_), .C(_12812_), .Y(_12814_) );
	AOI21X1 AOI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_11606_), .B(_12810_), .C(_12814_), .Y(_12815_) );
	NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(_12809_), .B(_12815_), .C(_12804_), .Y(_12816_) );
	INVX1 INVX1_2035 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .Y(_12817_) );
	NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_11606_), .Y(_12818_) );
	NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_11612_), .Y(_12819_) );
	NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_12818_), .B(_12819_), .Y(_12820_) );
	AOI21X1 AOI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_12784_), .B(_12817_), .C(_12820_), .Y(_12821_) );
	NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12820_), .C(_12784_), .Y(_12822_) );
	NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf0), .B(_12822_), .Y(_12823_) );
	OAI21X1 OAI21X1_5224 ( .gnd(gnd), .vdd(vdd), .A(_12821_), .B(_12823_), .C(_13398__bF_buf5), .Y(_12824_) );
	OAI21X1 OAI21X1_5225 ( .gnd(gnd), .vdd(vdd), .A(_12769_), .B(_13391__bF_buf4), .C(_13441__bF_buf1), .Y(_12825_) );
	OAI21X1 OAI21X1_5226 ( .gnd(gnd), .vdd(vdd), .A(_12824_), .B(_12816_), .C(_12825_), .Y(_12826_) );
	AOI21X1 AOI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_12826_), .B(_12803_), .C(rst_bF_buf64), .Y(_11292__17_) );
	INVX2 INVX2_175 ( .gnd(gnd), .vdd(vdd), .A(data_rd_19_), .Y(_12827_) );
	MUX2X1 MUX2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(_12800_), .S(_13416__bF_buf3), .Y(_12828_) );
	AOI21X1 AOI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_12769_), .B(_13415__bF_buf5), .C(_13392__bF_buf6), .Y(_12829_) );
	OAI21X1 OAI21X1_5227 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf4), .B(_12828_), .C(_12829_), .Y(_12830_) );
	OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_12783_), .B(_12820_), .Y(_12831_) );
	INVX1 INVX1_2036 ( .gnd(gnd), .vdd(vdd), .A(_12818_), .Y(_12832_) );
	AOI21X1 AOI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_12819_), .C(_12832_), .Y(_12833_) );
	OAI21X1 OAI21X1_5228 ( .gnd(gnd), .vdd(vdd), .A(_12831_), .B(_12779_), .C(_12833_), .Y(_12834_) );
	INVX1 INVX1_2037 ( .gnd(gnd), .vdd(vdd), .A(_12834_), .Y(_12835_) );
	NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_11662_), .Y(_12836_) );
	NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_11633_), .Y(_12837_) );
	NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_12837_), .B(_12836_), .Y(_12838_) );
	AOI21X1 AOI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_12835_), .B(_12838_), .C(_12294_), .Y(_12839_) );
	OAI21X1 OAI21X1_5229 ( .gnd(gnd), .vdd(vdd), .A(_12835_), .B(_12838_), .C(_12839_), .Y(_12840_) );
	OAI21X1 OAI21X1_5230 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf2), .B(addp_bF_buf2), .C(_11646_), .Y(_12841_) );
	AOI21X1 AOI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_12297__bF_buf3), .C(_12630_), .Y(_12842_) );
	OAI21X1 OAI21X1_5231 ( .gnd(gnd), .vdd(vdd), .A(_13458__bF_buf0), .B(_13466__bF_buf2), .C(biu_biu_data_out_18_), .Y(_12843_) );
	AOI21X1 AOI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_12333_), .C(_12626_), .Y(_12844_) );
	OAI21X1 OAI21X1_5232 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .B(_11662_), .C(_12290__bF_buf3), .Y(_12845_) );
	AOI22X1 AOI22X1_675 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_18_), .C(csr_18_), .D(_12305__bF_buf1), .Y(_12846_) );
	NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(_12843_), .B(_12846_), .C(_12845_), .Y(_12847_) );
	AOI21X1 AOI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_11662_), .B(_12842_), .C(_12847_), .Y(_12848_) );
	NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(_12840_), .B(_12848_), .C(_12841_), .Y(_12849_) );
	NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(_12807_), .Y(_12850_) );
	NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .B(biu_pc_18_), .C(_12805_), .Y(_12851_) );
	OAI21X1 OAI21X1_5233 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_ins_dec_jal_bF_buf5), .C(_12851_), .Y(_12852_) );
	OAI21X1 OAI21X1_5234 ( .gnd(gnd), .vdd(vdd), .A(_12850_), .B(_12852_), .C(_13398__bF_buf4), .Y(_12853_) );
	OAI21X1 OAI21X1_5235 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_13391__bF_buf3), .C(_13441__bF_buf0), .Y(_12854_) );
	OAI21X1 OAI21X1_5236 ( .gnd(gnd), .vdd(vdd), .A(_12853_), .B(_12849_), .C(_12854_), .Y(_12855_) );
	AOI21X1 AOI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_12855_), .B(_12830_), .C(rst_bF_buf63), .Y(_11292__18_) );
	INVX2 INVX2_176 ( .gnd(gnd), .vdd(vdd), .A(data_rd_20_), .Y(_12856_) );
	MUX2X1 MUX2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_12856_), .B(_12827_), .S(_13416__bF_buf2), .Y(_12857_) );
	AOI21X1 AOI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_13415__bF_buf3), .C(_13392__bF_buf5), .Y(_12858_) );
	OAI21X1 OAI21X1_5237 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf2), .B(_12857_), .C(_12858_), .Y(_12859_) );
	OAI21X1 OAI21X1_5238 ( .gnd(gnd), .vdd(vdd), .A(_12838_), .B(_12835_), .C(_12836_), .Y(_12860_) );
	NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_11666_), .Y(_12861_) );
	NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_12223_), .Y(_12862_) );
	OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_12861_), .B(_12862_), .Y(_12863_) );
	INVX1 INVX1_2038 ( .gnd(gnd), .vdd(vdd), .A(_12863_), .Y(_12864_) );
	OAI21X1 OAI21X1_5239 ( .gnd(gnd), .vdd(vdd), .A(_12864_), .B(_12860_), .C(csr_gpr_iu_ins_dec_subp_bF_buf3), .Y(_12865_) );
	AOI21X1 AOI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_12860_), .B(_12864_), .C(_12865_), .Y(_12866_) );
	OAI21X1 OAI21X1_5240 ( .gnd(gnd), .vdd(vdd), .A(_11667_), .B(_12851_), .C(_12337__bF_buf2), .Y(_12867_) );
	AOI21X1 AOI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_11667_), .B(_12851_), .C(_12867_), .Y(_12868_) );
	OAI21X1 OAI21X1_5241 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_12291__bF_buf0), .C(_12757_), .Y(_12869_) );
	OAI21X1 OAI21X1_5242 ( .gnd(gnd), .vdd(vdd), .A(_12869_), .B(_12223_), .C(_12290__bF_buf2), .Y(_12870_) );
	AOI21X1 AOI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_12297__bF_buf2), .C(_12630_), .Y(_12871_) );
	NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(csr_19_), .B(_12305__bF_buf0), .Y(_12872_) );
	AOI21X1 AOI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_19_), .C(_13695__bF_buf3), .Y(_12873_) );
	NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(_12222_), .B(_12872_), .C(_12873_), .Y(_12874_) );
	AOI21X1 AOI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_12223_), .B(_12871_), .C(_12874_), .Y(_12875_) );
	NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_12870_), .B(_12875_), .Y(_12876_) );
	NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_12876_), .B(_12868_), .Y(_12877_) );
	OAI21X1 OAI21X1_5243 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11673_), .C(_12877_), .Y(_12878_) );
	OAI21X1 OAI21X1_5244 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(_13391__bF_buf2), .C(_13441__bF_buf4), .Y(_12879_) );
	OAI21X1 OAI21X1_5245 ( .gnd(gnd), .vdd(vdd), .A(_12866_), .B(_12878_), .C(_12879_), .Y(_12880_) );
	AOI21X1 AOI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12859_), .C(rst_bF_buf62), .Y(_11292__19_) );
	INVX2 INVX2_177 ( .gnd(gnd), .vdd(vdd), .A(data_rd_21_), .Y(_12881_) );
	MUX2X1 MUX2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12856_), .S(_13416__bF_buf1), .Y(_12882_) );
	AOI21X1 AOI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(_13415__bF_buf1), .C(_13392__bF_buf4), .Y(_12883_) );
	OAI21X1 OAI21X1_5246 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf0), .B(_12882_), .C(_12883_), .Y(_12884_) );
	OAI21X1 OAI21X1_5247 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_19_), .B(_11666_), .C(_12836_), .Y(_12885_) );
	OAI21X1 OAI21X1_5248 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_12223_), .C(_12885_), .Y(_12886_) );
	OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_12863_), .B(_12838_), .Y(_12887_) );
	OAI21X1 OAI21X1_5249 ( .gnd(gnd), .vdd(vdd), .A(_12833_), .B(_12887_), .C(_12886_), .Y(_12888_) );
	INVX1 INVX1_2039 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .Y(_12889_) );
	NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_12887_), .B(_12831_), .Y(_12890_) );
	INVX1 INVX1_2040 ( .gnd(gnd), .vdd(vdd), .A(_12890_), .Y(_12891_) );
	OAI21X1 OAI21X1_5250 ( .gnd(gnd), .vdd(vdd), .A(_12891_), .B(_12779_), .C(_12889_), .Y(_12892_) );
	NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_11698_), .Y(_12893_) );
	NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(_11699_), .Y(_12894_) );
	AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_12894_), .B(_12893_), .Y(_12895_) );
	AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_12892_), .B(_12895_), .Y(_12896_) );
	OAI21X1 OAI21X1_5251 ( .gnd(gnd), .vdd(vdd), .A(_12895_), .B(_12892_), .C(csr_gpr_iu_ins_dec_subp_bF_buf2), .Y(_12897_) );
	OAI21X1 OAI21X1_5252 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf1), .B(addp_bF_buf1), .C(_11706_), .Y(_12898_) );
	AOI21X1 AOI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_12297__bF_buf1), .C(_12630_), .Y(_12899_) );
	AOI21X1 AOI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_12333_), .C(_12626_), .Y(_12900_) );
	OAI21X1 OAI21X1_5253 ( .gnd(gnd), .vdd(vdd), .A(_12900_), .B(_11698_), .C(_12290__bF_buf1), .Y(_12901_) );
	AOI22X1 AOI22X1_676 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_20_bF_buf3), .C(csr_20_), .D(_12305__bF_buf4), .Y(_12902_) );
	NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(_11697_), .B(_12902_), .C(_12901_), .Y(_12903_) );
	AOI21X1 AOI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .B(_12899_), .C(_12903_), .Y(_12904_) );
	AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .B(_12904_), .Y(_12905_) );
	OAI21X1 OAI21X1_5254 ( .gnd(gnd), .vdd(vdd), .A(_12896_), .B(_12897_), .C(_12905_), .Y(_12906_) );
	INVX1 INVX1_2041 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .Y(_12907_) );
	NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_11667_), .B(_12907_), .C(_12851_), .Y(_12908_) );
	NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .B(biu_pc_19_), .C(_12807_), .Y(_12909_) );
	INVX1 INVX1_2042 ( .gnd(gnd), .vdd(vdd), .A(_12909_), .Y(_12910_) );
	OAI21X1 OAI21X1_5255 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .B(_12910_), .C(_12337__bF_buf1), .Y(_12911_) );
	OAI21X1 OAI21X1_5256 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .B(_12911_), .C(_13398__bF_buf3), .Y(_12912_) );
	OAI21X1 OAI21X1_5257 ( .gnd(gnd), .vdd(vdd), .A(_12856_), .B(_13391__bF_buf1), .C(_13441__bF_buf3), .Y(_12913_) );
	OAI21X1 OAI21X1_5258 ( .gnd(gnd), .vdd(vdd), .A(_12912_), .B(_12906_), .C(_12913_), .Y(_12914_) );
	AOI21X1 AOI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_12914_), .B(_12884_), .C(rst_bF_buf61), .Y(_11292__20_) );
	INVX2 INVX2_178 ( .gnd(gnd), .vdd(vdd), .A(data_rd_22_), .Y(_12915_) );
	MUX2X1 MUX2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_12881_), .S(_13416__bF_buf0), .Y(_12916_) );
	AOI21X1 AOI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_12856_), .B(_13415__bF_buf6), .C(_13392__bF_buf3), .Y(_12917_) );
	OAI21X1 OAI21X1_5259 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf5), .B(_12916_), .C(_12917_), .Y(_12918_) );
	INVX1 INVX1_2043 ( .gnd(gnd), .vdd(vdd), .A(_12893_), .Y(_12919_) );
	NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_12919_), .B(_12896_), .Y(_12920_) );
	NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_11732_), .Y(_12921_) );
	INVX1 INVX1_2044 ( .gnd(gnd), .vdd(vdd), .A(_12921_), .Y(_12922_) );
	NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(_11732_), .Y(_12923_) );
	AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .B(_12923_), .Y(_12924_) );
	INVX1 INVX1_2045 ( .gnd(gnd), .vdd(vdd), .A(_12924_), .Y(_12925_) );
	AOI21X1 AOI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_12920_), .B(_12925_), .C(_12294_), .Y(_12926_) );
	OAI21X1 OAI21X1_5260 ( .gnd(gnd), .vdd(vdd), .A(_12920_), .B(_12925_), .C(_12926_), .Y(_12927_) );
	OAI21X1 OAI21X1_5261 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf0), .B(addp_bF_buf0), .C(_11736_), .Y(_12928_) );
	AOI21X1 AOI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_12297__bF_buf0), .C(_12630_), .Y(_12929_) );
	OAI21X1 OAI21X1_5262 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_12291__bF_buf3), .C(_12757_), .Y(_12930_) );
	OAI21X1 OAI21X1_5263 ( .gnd(gnd), .vdd(vdd), .A(_12930_), .B(_11726_), .C(_12290__bF_buf0), .Y(_12931_) );
	AOI22X1 AOI22X1_677 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_21_bF_buf3), .C(csr_21_), .D(_12305__bF_buf3), .Y(_12932_) );
	NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_12932_), .C(_12931_), .Y(_12933_) );
	AOI21X1 AOI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_12929_), .C(_12933_), .Y(_12934_) );
	NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(_12927_), .B(_12934_), .C(_12928_), .Y(_12935_) );
	INVX1 INVX1_2046 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .Y(_12936_) );
	NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_12907_), .B(_12936_), .C(_12909_), .Y(_12937_) );
	NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12937_), .Y(_12938_) );
	OAI21X1 OAI21X1_5264 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .B(_12908_), .C(_12938_), .Y(_12939_) );
	NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf2), .B(_12939_), .Y(_12940_) );
	OAI21X1 OAI21X1_5265 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_13391__bF_buf0), .C(_13441__bF_buf2), .Y(_12941_) );
	OAI21X1 OAI21X1_5266 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .B(_12935_), .C(_12941_), .Y(_12942_) );
	AOI21X1 AOI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_12942_), .B(_12918_), .C(rst_bF_buf60), .Y(_11292__21_) );
	INVX2 INVX2_179 ( .gnd(gnd), .vdd(vdd), .A(data_rd_23_), .Y(_12943_) );
	MUX2X1 MUX2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_12915_), .S(_13416__bF_buf4), .Y(_12944_) );
	AOI21X1 AOI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_13415__bF_buf4), .C(_13392__bF_buf2), .Y(_12945_) );
	OAI21X1 OAI21X1_5267 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf3), .B(_12944_), .C(_12945_), .Y(_12946_) );
	AOI21X1 AOI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_11768_), .B(_11767_), .C(_12348_), .Y(_12947_) );
	OAI21X1 OAI21X1_5268 ( .gnd(gnd), .vdd(vdd), .A(_12921_), .B(_12919_), .C(_12923_), .Y(_12948_) );
	INVX1 INVX1_2047 ( .gnd(gnd), .vdd(vdd), .A(_12948_), .Y(_12949_) );
	NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_12895_), .B(_12924_), .Y(_12950_) );
	INVX1 INVX1_2048 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .Y(_12951_) );
	AOI21X1 AOI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_12892_), .B(_12951_), .C(_12949_), .Y(_12952_) );
	NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_11753_), .Y(_12953_) );
	INVX1 INVX1_2049 ( .gnd(gnd), .vdd(vdd), .A(_12953_), .Y(_12954_) );
	NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_11753_), .Y(_12955_) );
	AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_12954_), .B(_12955_), .Y(_12956_) );
	INVX1 INVX1_2050 ( .gnd(gnd), .vdd(vdd), .A(_12956_), .Y(_12957_) );
	AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_12952_), .B(_12957_), .Y(_12958_) );
	OAI21X1 OAI21X1_5269 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .B(_12952_), .C(csr_gpr_iu_ins_dec_subp_bF_buf1), .Y(_12959_) );
	OAI21X1 OAI21X1_5270 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_12937_), .C(_12337__bF_buf0), .Y(_12960_) );
	AOI21X1 AOI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(_12937_), .C(_12960_), .Y(_12961_) );
	OAI21X1 OAI21X1_5271 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .B(_12291__bF_buf2), .C(_12757_), .Y(_12962_) );
	OAI21X1 OAI21X1_5272 ( .gnd(gnd), .vdd(vdd), .A(_12962_), .B(_11759_), .C(_12290__bF_buf4), .Y(_12963_) );
	AOI21X1 AOI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .B(_12297__bF_buf4), .C(_12630_), .Y(_12964_) );
	NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(csr_22_), .B(_12305__bF_buf2), .Y(_12965_) );
	AOI21X1 AOI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_22_bF_buf1), .C(_13695__bF_buf2), .Y(_12966_) );
	NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(_11758_), .B(_12965_), .C(_12966_), .Y(_12967_) );
	AOI21X1 AOI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_12964_), .C(_12967_), .Y(_12968_) );
	NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_12963_), .B(_12968_), .Y(_12969_) );
	NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_12969_), .B(_12961_), .Y(_12970_) );
	OAI21X1 OAI21X1_5273 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .B(_12959_), .C(_12970_), .Y(_12971_) );
	OAI21X1 OAI21X1_5274 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_13391__bF_buf7), .C(_13441__bF_buf1), .Y(_12972_) );
	OAI21X1 OAI21X1_5275 ( .gnd(gnd), .vdd(vdd), .A(_12971_), .B(_12947_), .C(_12972_), .Y(_12973_) );
	AOI21X1 AOI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_12973_), .B(_12946_), .C(rst_bF_buf59), .Y(_11292__22_) );
	INVX2 INVX2_180 ( .gnd(gnd), .vdd(vdd), .A(data_rd_24_), .Y(_12974_) );
	MUX2X1 MUX2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12943_), .S(_13416__bF_buf3), .Y(_12975_) );
	AOI21X1 AOI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_13415__bF_buf2), .C(_13392__bF_buf1), .Y(_12976_) );
	OAI21X1 OAI21X1_5276 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf1), .B(_12975_), .C(_12976_), .Y(_12977_) );
	OAI21X1 OAI21X1_5277 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .B(_12952_), .C(_12954_), .Y(_12978_) );
	NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_23_), .B(_11793_), .Y(_12979_) );
	NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_11799_), .Y(_12980_) );
	NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_12979_), .B(_12980_), .Y(_12981_) );
	AOI21X1 AOI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_12981_), .C(_12294_), .Y(_12982_) );
	OAI21X1 OAI21X1_5278 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_12981_), .C(_12982_), .Y(_12983_) );
	NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(_11806_), .B(_12405_), .C(_11804_), .Y(_12984_) );
	AOI21X1 AOI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_12297__bF_buf3), .C(_12630_), .Y(_12985_) );
	OAI21X1 OAI21X1_5279 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_12291__bF_buf1), .C(_12757_), .Y(_12986_) );
	OAI21X1 OAI21X1_5280 ( .gnd(gnd), .vdd(vdd), .A(_12986_), .B(_11799_), .C(_12290__bF_buf3), .Y(_12987_) );
	AOI22X1 AOI22X1_678 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_23_), .C(csr_23_), .D(_12305__bF_buf1), .Y(_12988_) );
	NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .B(_12988_), .C(_12987_), .Y(_12989_) );
	AOI21X1 AOI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_12985_), .C(_12989_), .Y(_12990_) );
	NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(_12983_), .B(_12990_), .C(_12984_), .Y(_12991_) );
	INVX1 INVX1_2051 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .Y(_12992_) );
	NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .B(biu_pc_22_), .C(_12908_), .Y(_12993_) );
	AOI21X1 AOI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_12993_), .B(_12992_), .C(_12306_), .Y(_12994_) );
	OAI21X1 OAI21X1_5281 ( .gnd(gnd), .vdd(vdd), .A(_12992_), .B(_12993_), .C(_12994_), .Y(_12995_) );
	NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_13398__bF_buf1), .B(_12995_), .Y(_12996_) );
	OAI21X1 OAI21X1_5282 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_13391__bF_buf6), .C(_13441__bF_buf0), .Y(_12997_) );
	OAI21X1 OAI21X1_5283 ( .gnd(gnd), .vdd(vdd), .A(_12996_), .B(_12991_), .C(_12997_), .Y(_12998_) );
	AOI21X1 AOI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_12998_), .B(_12977_), .C(rst_bF_buf58), .Y(_11292__23_) );
	INVX2 INVX2_181 ( .gnd(gnd), .vdd(vdd), .A(data_rd_25_), .Y(_12999_) );
	MUX2X1 MUX2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_12999_), .B(_12974_), .S(_13416__bF_buf2), .Y(_13000_) );
	AOI21X1 AOI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_13415__bF_buf0), .C(_13392__bF_buf0), .Y(_13001_) );
	OAI21X1 OAI21X1_5284 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf6), .B(_13000_), .C(_13001_), .Y(_13002_) );
	NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_12981_), .B(_12956_), .Y(_13003_) );
	NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_13003_), .Y(_13004_) );
	NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_13004_), .B(_12890_), .Y(_13005_) );
	AOI21X1 AOI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_12981_), .B(_12953_), .C(_12979_), .Y(_13006_) );
	OAI21X1 OAI21X1_5285 ( .gnd(gnd), .vdd(vdd), .A(_12948_), .B(_13003_), .C(_13006_), .Y(_13007_) );
	AOI21X1 AOI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .B(_13004_), .C(_13007_), .Y(_13008_) );
	OAI21X1 OAI21X1_5286 ( .gnd(gnd), .vdd(vdd), .A(_13005_), .B(_12779_), .C(_13008_), .Y(_13009_) );
	XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(csr_gpr_iu_rs2_24_), .Y(_13010_) );
	OAI21X1 OAI21X1_5287 ( .gnd(gnd), .vdd(vdd), .A(_13010_), .B(_13009_), .C(csr_gpr_iu_ins_dec_subp_bF_buf0), .Y(_13011_) );
	AOI21X1 AOI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .B(_13010_), .C(_13011_), .Y(_13012_) );
	INVX1 INVX1_2052 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .Y(_13013_) );
	INVX2 INVX2_182 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .Y(_13014_) );
	NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_12992_), .B(_13014_), .C(_12993_), .Y(_13015_) );
	INVX1 INVX1_2053 ( .gnd(gnd), .vdd(vdd), .A(_13015_), .Y(_13016_) );
	NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .B(biu_pc_23_), .C(_12937_), .Y(_13017_) );
	AOI21X1 AOI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_13017_), .B(_13014_), .C(_12306_), .Y(_13018_) );
	AOI21X1 AOI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_12297__bF_buf2), .C(_12630_), .Y(_13019_) );
	OAI21X1 OAI21X1_5288 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf2), .B(_13019_), .C(_11834_), .Y(_13020_) );
	OAI21X1 OAI21X1_5289 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .B(_12291__bF_buf0), .C(_12698_), .Y(_13021_) );
	NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(csr_24_), .B(_12305__bF_buf0), .Y(_13022_) );
	AOI21X1 AOI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_24_), .C(_13695__bF_buf1), .Y(_13023_) );
	NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(_13021_), .B(_13022_), .C(_13023_), .Y(_13024_) );
	INVX1 INVX1_2054 ( .gnd(gnd), .vdd(vdd), .A(_13024_), .Y(_13025_) );
	NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_13020_), .C(_13025_), .Y(_13026_) );
	AOI21X1 AOI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_13018_), .C(_13026_), .Y(_13027_) );
	OAI21X1 OAI21X1_5290 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_13013_), .C(_13027_), .Y(_13028_) );
	OAI21X1 OAI21X1_5291 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_13391__bF_buf5), .C(_13441__bF_buf4), .Y(_13029_) );
	OAI21X1 OAI21X1_5292 ( .gnd(gnd), .vdd(vdd), .A(_13012_), .B(_13028_), .C(_13029_), .Y(_13030_) );
	AOI21X1 AOI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_13030_), .B(_13002_), .C(rst_bF_buf57), .Y(_11292__24_) );
	INVX2 INVX2_183 ( .gnd(gnd), .vdd(vdd), .A(data_rd_26_), .Y(_13031_) );
	MUX2X1 MUX2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .B(_12999_), .S(_13416__bF_buf1), .Y(_13032_) );
	AOI21X1 AOI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_13415__bF_buf5), .C(_13392__bF_buf7), .Y(_13033_) );
	OAI21X1 OAI21X1_5293 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf4), .B(_13032_), .C(_13033_), .Y(_13034_) );
	OAI21X1 OAI21X1_5294 ( .gnd(gnd), .vdd(vdd), .A(_12999_), .B(_13391__bF_buf4), .C(_13441__bF_buf3), .Y(_13035_) );
	NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11867_), .Y(_13036_) );
	NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_11860_), .Y(_13037_) );
	NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_11871_), .Y(_13038_) );
	NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .B(_13038_), .Y(_13039_) );
	INVX1 INVX1_2055 ( .gnd(gnd), .vdd(vdd), .A(_13039_), .Y(_13040_) );
	NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_13010_), .B(_13009_), .Y(_13041_) );
	OAI21X1 OAI21X1_5295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .B(_11842_), .C(_13041_), .Y(_13042_) );
	XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_13042_), .B(_13040_), .Y(_13043_) );
	INVX1 INVX1_2056 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .Y(_13044_) );
	NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_13014_), .B(_13044_), .C(_13017_), .Y(_13045_) );
	NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_13045_), .Y(_13046_) );
	OAI21X1 OAI21X1_5296 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .B(_13015_), .C(_13046_), .Y(_13047_) );
	OAI21X1 OAI21X1_5297 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .B(_12291__bF_buf3), .C(_12757_), .Y(_13048_) );
	OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(_13048_), .Y(_13049_) );
	OAI21X1 OAI21X1_5298 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_12296_), .C(_12631_), .Y(_13050_) );
	INVX2 INVX2_184 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .Y(_13051_) );
	INVX1 INVX1_2057 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf0), .Y(_13052_) );
	OAI21X1 OAI21X1_5299 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13052_), .C(_13398__bF_buf0), .Y(_13053_) );
	AOI21X1 AOI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(csr_25_), .B(_12305__bF_buf4), .C(_13053_), .Y(_13054_) );
	AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_13054_), .B(_11859_), .Y(_13055_) );
	OAI21X1 OAI21X1_5300 ( .gnd(gnd), .vdd(vdd), .A(_11871_), .B(_13050_), .C(_13055_), .Y(_13056_) );
	AOI21X1 AOI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf1), .B(_13049_), .C(_13056_), .Y(_13057_) );
	AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(_13047_), .B(_13057_), .Y(_13058_) );
	OAI21X1 OAI21X1_5301 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_13043_), .C(_13058_), .Y(_13059_) );
	OAI21X1 OAI21X1_5302 ( .gnd(gnd), .vdd(vdd), .A(_13036_), .B(_13059_), .C(_13035_), .Y(_13060_) );
	AOI21X1 AOI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_13060_), .B(_13034_), .C(rst_bF_buf56), .Y(_11292__25_) );
	INVX2 INVX2_185 ( .gnd(gnd), .vdd(vdd), .A(data_rd_27_), .Y(_13061_) );
	MUX2X1 MUX2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13031_), .S(_13416__bF_buf0), .Y(_13062_) );
	AOI21X1 AOI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_12999_), .B(_13415__bF_buf3), .C(_13392__bF_buf6), .Y(_13063_) );
	OAI21X1 OAI21X1_5303 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf2), .B(_13062_), .C(_13063_), .Y(_13064_) );
	OAI21X1 OAI21X1_5304 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(_13045_), .C(_12337__bF_buf3), .Y(_13065_) );
	AOI21X1 AOI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(_13045_), .C(_13065_), .Y(_13066_) );
	OAI21X1 OAI21X1_5305 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_12291__bF_buf2), .C(_12757_), .Y(_13067_) );
	OAI21X1 OAI21X1_5306 ( .gnd(gnd), .vdd(vdd), .A(_13067_), .B(_11886_), .C(_12290__bF_buf0), .Y(_13068_) );
	AOI21X1 AOI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_12297__bF_buf1), .C(_12630_), .Y(_13069_) );
	NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(csr_26_), .B(_12305__bF_buf3), .Y(_13070_) );
	NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_26_bF_buf2), .Y(_13071_) );
	NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(_13070_), .B(_13071_), .C(_11885_), .Y(_13072_) );
	AOI21X1 AOI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_11886_), .B(_13069_), .C(_13072_), .Y(_13073_) );
	NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_13068_), .B(_13073_), .Y(_13074_) );
	NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_13074_), .B(_13066_), .Y(_13075_) );
	OAI21X1 OAI21X1_5307 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_11900_), .C(_13075_), .Y(_13076_) );
	NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_13010_), .B(_13040_), .Y(_13077_) );
	INVX1 INVX1_2058 ( .gnd(gnd), .vdd(vdd), .A(_13077_), .Y(_13078_) );
	NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_11834_), .Y(_13079_) );
	OAI21X1 OAI21X1_5308 ( .gnd(gnd), .vdd(vdd), .A(_13079_), .B(_13039_), .C(_13037_), .Y(_13080_) );
	AOI21X1 AOI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .B(_13078_), .C(_13080_), .Y(_13081_) );
	NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_11886_), .Y(_13082_) );
	NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_11904_), .Y(_13083_) );
	NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_13082_), .B(_13083_), .Y(_13084_) );
	AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_13081_), .B(_13084_), .Y(_13085_) );
	OAI21X1 OAI21X1_5309 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_13081_), .C(csr_gpr_iu_ins_dec_subp_bF_buf3), .Y(_13086_) );
	OAI21X1 OAI21X1_5310 ( .gnd(gnd), .vdd(vdd), .A(_13085_), .B(_13086_), .C(_13398__bF_buf6), .Y(_13087_) );
	OAI21X1 OAI21X1_5311 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .B(_13391__bF_buf3), .C(_13441__bF_buf2), .Y(_13088_) );
	OAI21X1 OAI21X1_5312 ( .gnd(gnd), .vdd(vdd), .A(_13087_), .B(_13076_), .C(_13088_), .Y(_13089_) );
	AOI21X1 AOI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_13089_), .B(_13064_), .C(rst_bF_buf55), .Y(_11292__26_) );
	INVX2 INVX2_186 ( .gnd(gnd), .vdd(vdd), .A(data_rd_28_), .Y(_13090_) );
	MUX2X1 MUX2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_13090_), .B(_13061_), .S(_13416__bF_buf4), .Y(_13091_) );
	AOI21X1 AOI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .B(_13415__bF_buf1), .C(_13392__bF_buf5), .Y(_13092_) );
	OAI21X1 OAI21X1_5313 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf0), .B(_13091_), .C(_13092_), .Y(_13093_) );
	OAI21X1 OAI21X1_5314 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13391__bF_buf2), .C(_13441__bF_buf1), .Y(_13094_) );
	AOI21X1 AOI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_11927_), .B(_11928_), .C(_12348_), .Y(_13095_) );
	OAI21X1 OAI21X1_5315 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_13081_), .C(_13082_), .Y(_13096_) );
	XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_13508_), .Y(_13097_) );
	AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_13096_), .B(_13097_), .Y(_13098_) );
	OAI21X1 OAI21X1_5316 ( .gnd(gnd), .vdd(vdd), .A(_13097_), .B(_13096_), .C(csr_gpr_iu_ins_dec_subp_bF_buf2), .Y(_13099_) );
	NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .B(biu_pc_27_), .C(_13045_), .Y(_13100_) );
	INVX1 INVX1_2059 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .Y(_13101_) );
	NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .B(biu_pc_26_), .C(_13015_), .Y(_13102_) );
	AOI21X1 AOI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_13102_), .B(_13101_), .C(_12306_), .Y(_13103_) );
	OAI21X1 OAI21X1_5317 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_12291__bF_buf1), .C(_12757_), .Y(_13104_) );
	OAI21X1 OAI21X1_5318 ( .gnd(gnd), .vdd(vdd), .A(_13104_), .B(_11921_), .C(_12290__bF_buf4), .Y(_13105_) );
	AOI21X1 AOI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_12297__bF_buf0), .C(_12630_), .Y(_13106_) );
	NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(csr_27_), .B(_12305__bF_buf2), .Y(_13107_) );
	AOI21X1 AOI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lui), .B(biu_ins_27_bF_buf1), .C(_13695__bF_buf0), .Y(_13108_) );
	NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(_11920_), .B(_13107_), .C(_13108_), .Y(_13109_) );
	AOI21X1 AOI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .B(_13106_), .C(_13109_), .Y(_13110_) );
	NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_13105_), .B(_13110_), .Y(_13111_) );
	AOI21X1 AOI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_13103_), .B(_13100_), .C(_13111_), .Y(_13112_) );
	OAI21X1 OAI21X1_5319 ( .gnd(gnd), .vdd(vdd), .A(_13098_), .B(_13099_), .C(_13112_), .Y(_13113_) );
	OAI21X1 OAI21X1_5320 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13095_), .C(_13094_), .Y(_13114_) );
	AOI21X1 AOI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_13114_), .B(_13093_), .C(rst_bF_buf54), .Y(_11292__27_) );
	INVX2 INVX2_187 ( .gnd(gnd), .vdd(vdd), .A(data_rd_29_), .Y(_13115_) );
	MUX2X1 MUX2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13090_), .S(_13416__bF_buf3), .Y(_13116_) );
	AOI21X1 AOI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13415__bF_buf6), .C(_13392__bF_buf4), .Y(_13117_) );
	OAI21X1 OAI21X1_5321 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf5), .B(_13116_), .C(_13117_), .Y(_13118_) );
	INVX1 INVX1_2060 ( .gnd(gnd), .vdd(vdd), .A(_13100_), .Y(_13119_) );
	INVX1 INVX1_2061 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .Y(_13120_) );
	NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_13101_), .B(_13120_), .C(_13102_), .Y(_13121_) );
	NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_13121_), .Y(_13122_) );
	OAI21X1 OAI21X1_5322 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .B(_13119_), .C(_13122_), .Y(_13123_) );
	OAI21X1 OAI21X1_5323 ( .gnd(gnd), .vdd(vdd), .A(addi_bF_buf6), .B(addp_bF_buf4), .C(_11963_), .Y(_13124_) );
	OAI21X1 OAI21X1_5324 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_12291__bF_buf0), .C(_12757_), .Y(_13125_) );
	OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .B(_13125_), .Y(_13126_) );
	OAI21X1 OAI21X1_5325 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_12296_), .C(_12631_), .Y(_13127_) );
	INVX1 INVX1_2062 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf2), .Y(_13128_) );
	OAI21X1 OAI21X1_5326 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13128_), .C(_11952_), .Y(_13129_) );
	AOI21X1 AOI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(csr_28_), .B(_12305__bF_buf1), .C(_13129_), .Y(_13130_) );
	OAI21X1 OAI21X1_5327 ( .gnd(gnd), .vdd(vdd), .A(_13127_), .B(_11954_), .C(_13130_), .Y(_13131_) );
	AOI21X1 AOI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf3), .B(_13126_), .C(_13131_), .Y(_13132_) );
	NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(_13124_), .B(_13132_), .C(_13123_), .Y(_13133_) );
	NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(_13082_), .B(_13083_), .C(_13097_), .Y(_13134_) );
	NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(_13077_), .Y(_13135_) );
	INVX1 INVX1_2063 ( .gnd(gnd), .vdd(vdd), .A(_13080_), .Y(_13136_) );
	OAI21X1 OAI21X1_5328 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_27_), .B(_11932_), .C(_13082_), .Y(_13137_) );
	OAI21X1 OAI21X1_5329 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_11921_), .C(_13137_), .Y(_13138_) );
	OAI21X1 OAI21X1_5330 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(_13136_), .C(_13138_), .Y(_13139_) );
	AOI21X1 AOI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .B(_13135_), .C(_13139_), .Y(_13140_) );
	NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_11954_), .Y(_13141_) );
	NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_11953_), .Y(_13142_) );
	NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_13142_), .B(_13141_), .Y(_13143_) );
	INVX1 INVX1_2064 ( .gnd(gnd), .vdd(vdd), .A(_13143_), .Y(_13144_) );
	NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_13144_), .B(_13140_), .Y(_13145_) );
	OAI21X1 OAI21X1_5331 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13142_), .C(_13140_), .Y(_13146_) );
	NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_subp_bF_buf1), .B(_13146_), .Y(_13147_) );
	OAI21X1 OAI21X1_5332 ( .gnd(gnd), .vdd(vdd), .A(_13145_), .B(_13147_), .C(_13398__bF_buf5), .Y(_13148_) );
	OAI21X1 OAI21X1_5333 ( .gnd(gnd), .vdd(vdd), .A(_13090_), .B(_13391__bF_buf1), .C(_13441__bF_buf0), .Y(_13149_) );
	OAI21X1 OAI21X1_5334 ( .gnd(gnd), .vdd(vdd), .A(_13148_), .B(_13133_), .C(_13149_), .Y(_13150_) );
	AOI21X1 AOI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_13150_), .B(_13118_), .C(rst_bF_buf53), .Y(_11292__28_) );
	INVX2 INVX2_188 ( .gnd(gnd), .vdd(vdd), .A(data_rd_30_), .Y(_13151_) );
	MUX2X1 MUX2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13115_), .S(_13416__bF_buf2), .Y(_13152_) );
	AOI21X1 AOI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_13090_), .B(_13415__bF_buf4), .C(_13392__bF_buf3), .Y(_13153_) );
	OAI21X1 OAI21X1_5335 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf3), .B(_13152_), .C(_13153_), .Y(_13154_) );
	NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .B(_11984_), .Y(_13155_) );
	NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_11983_), .Y(_13156_) );
	NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_13156_), .B(_13155_), .Y(_13157_) );
	INVX1 INVX1_2065 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .Y(_13158_) );
	OAI21X1 OAI21X1_5336 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13145_), .C(_13158_), .Y(_13159_) );
	NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13145_), .Y(_13160_) );
	NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .B(_13160_), .Y(_13161_) );
	AOI21X1 AOI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_13161_), .B(_13159_), .C(_12294_), .Y(_13162_) );
	NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(_11994_), .B(_12405_), .C(_11993_), .Y(_13163_) );
	INVX1 INVX1_2066 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .Y(_13164_) );
	NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_13120_), .B(_13164_), .C(_13100_), .Y(_13165_) );
	OAI21X1 OAI21X1_5337 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(_13121_), .C(_12337__bF_buf2), .Y(_13166_) );
	OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13165_), .Y(_13167_) );
	OAI21X1 OAI21X1_5338 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_12291__bF_buf3), .C(_12757_), .Y(_13168_) );
	OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_13168_), .Y(_13169_) );
	OAI21X1 OAI21X1_5339 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .B(_12296_), .C(_12631_), .Y(_13170_) );
	INVX1 INVX1_2067 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf3), .Y(_13171_) );
	OAI21X1 OAI21X1_5340 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13171_), .C(_13398__bF_buf4), .Y(_13172_) );
	AOI21X1 AOI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(csr_29_), .B(_12305__bF_buf0), .C(_13172_), .Y(_13173_) );
	AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_13173_), .B(_11982_), .Y(_13174_) );
	OAI21X1 OAI21X1_5341 ( .gnd(gnd), .vdd(vdd), .A(_11984_), .B(_13170_), .C(_13174_), .Y(_13175_) );
	AOI21X1 AOI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf2), .B(_13169_), .C(_13175_), .Y(_13176_) );
	NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(_13167_), .B(_13176_), .C(_13163_), .Y(_13177_) );
	OAI21X1 OAI21X1_5342 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13391__bF_buf0), .C(_13441__bF_buf4), .Y(_13178_) );
	OAI21X1 OAI21X1_5343 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .B(_13177_), .C(_13178_), .Y(_13179_) );
	AOI21X1 AOI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_13179_), .B(_13154_), .C(rst_bF_buf52), .Y(_11292__29_) );
	INVX1 INVX1_2068 ( .gnd(gnd), .vdd(vdd), .A(data_rd_31_), .Y(_13180_) );
	MUX2X1 MUX2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13151_), .S(_13416__bF_buf1), .Y(_13181_) );
	AOI21X1 AOI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13415__bF_buf2), .C(_13392__bF_buf2), .Y(_13182_) );
	OAI21X1 OAI21X1_5344 ( .gnd(gnd), .vdd(vdd), .A(_13415__bF_buf1), .B(_13181_), .C(_13182_), .Y(_13183_) );
	OAI21X1 OAI21X1_5345 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13391__bF_buf7), .C(_13441__bF_buf3), .Y(_13184_) );
	NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_13143_), .B(_13157_), .Y(_13185_) );
	AOI21X1 AOI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .B(_13141_), .C(_13155_), .Y(_13186_) );
	OAI21X1 OAI21X1_5346 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13140_), .C(_13186_), .Y(_13187_) );
	NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_12027_), .Y(_13188_) );
	NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_12017_), .Y(_13189_) );
	NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_13189_), .B(_13188_), .Y(_13190_) );
	XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_13187_), .B(_13190_), .Y(_13191_) );
	NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_13191_), .Y(_13192_) );
	AOI21X1 AOI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(biu_pc_30_), .C(_12306_), .Y(_13193_) );
	OAI21X1 OAI21X1_5347 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(_13165_), .C(_13193_), .Y(_13194_) );
	OAI21X1 OAI21X1_5348 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12021_), .C(_12405_), .Y(_13195_) );
	OAI21X1 OAI21X1_5349 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_12291__bF_buf2), .C(_12757_), .Y(_13196_) );
	OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_12017_), .B(_13196_), .Y(_13197_) );
	OAI21X1 OAI21X1_5350 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_12296_), .C(_12631_), .Y(_13198_) );
	INVX1 INVX1_2069 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf1), .Y(_13199_) );
	OAI21X1 OAI21X1_5351 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13199_), .C(_13398__bF_buf3), .Y(_13200_) );
	AOI21X1 AOI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(csr_30_), .B(_12305__bF_buf4), .C(_13200_), .Y(_13201_) );
	AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .B(_12016_), .Y(_13202_) );
	OAI21X1 OAI21X1_5352 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_13198_), .C(_13202_), .Y(_13203_) );
	AOI21X1 AOI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf1), .B(_13197_), .C(_13203_), .Y(_13204_) );
	NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(_13204_), .B(_13195_), .C(_13194_), .Y(_13205_) );
	OAI21X1 OAI21X1_5353 ( .gnd(gnd), .vdd(vdd), .A(_13192_), .B(_13205_), .C(_13184_), .Y(_13206_) );
	AOI21X1 AOI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_13206_), .B(_13183_), .C(rst_bF_buf51), .Y(_11292__30_) );
	OAI22X1 OAI22X1_824 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13414_), .C(_13180_), .D(_13418_), .Y(_13207_) );
	NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_13391__bF_buf6), .B(_13207_), .Y(_13208_) );
	AOI21X1 AOI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_13187_), .B(_13190_), .C(_13188_), .Y(_13209_) );
	XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .B(_13674_), .Y(_13210_) );
	OAI21X1 OAI21X1_5354 ( .gnd(gnd), .vdd(vdd), .A(_13210_), .B(_13209_), .C(csr_gpr_iu_ins_dec_subp_bF_buf0), .Y(_13211_) );
	AOI21X1 AOI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_13209_), .B(_13210_), .C(_13211_), .Y(_13212_) );
	NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(_12061_), .B(_12405_), .C(_12064_), .Y(_13213_) );
	NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(biu_pc_31_), .C(_13165_), .Y(_13214_) );
	INVX1 INVX1_2070 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .Y(_13215_) );
	NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(biu_pc_30_), .C(_13121_), .Y(_13216_) );
	NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_13215_), .B(_13216_), .Y(_13217_) );
	NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf1), .B(_13214_), .C(_13217_), .Y(_13218_) );
	OAI21X1 OAI21X1_5355 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_12291__bF_buf1), .C(_12757_), .Y(_13219_) );
	OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .B(_13219_), .Y(_13220_) );
	OAI21X1 OAI21X1_5356 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_12296_), .C(_12631_), .Y(_13221_) );
	INVX1 INVX1_2071 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .Y(_13222_) );
	OAI21X1 OAI21X1_5357 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13222_), .C(_13398__bF_buf2), .Y(_13223_) );
	AOI21X1 AOI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(csr_31_), .B(_12305__bF_buf3), .C(_13223_), .Y(_13224_) );
	AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .B(_12055_), .Y(_13225_) );
	OAI21X1 OAI21X1_5358 ( .gnd(gnd), .vdd(vdd), .A(_12068_), .B(_13221_), .C(_13225_), .Y(_13226_) );
	AOI21X1 AOI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_12290__bF_buf0), .B(_13220_), .C(_13226_), .Y(_13227_) );
	NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(_13227_), .B(_13218_), .C(_13213_), .Y(_13228_) );
	OAI21X1 OAI21X1_5359 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13391__bF_buf5), .C(_13441__bF_buf2), .Y(_13229_) );
	OAI21X1 OAI21X1_5360 ( .gnd(gnd), .vdd(vdd), .A(_13212_), .B(_13228_), .C(_13229_), .Y(_13230_) );
	AOI21X1 AOI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13208_), .C(rst_bF_buf50), .Y(_11292__31_) );
	NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_31_), .B(_12054_), .Y(_13231_) );
	NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_25_), .B(_11858_), .Y(_13232_) );
	NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_25_), .B(_13515_), .Y(_13233_) );
	NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_13232_), .B(_13233_), .Y(_13234_) );
	NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_24_), .B(_13516_), .Y(_13235_) );
	NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_24_), .B(_11832_), .Y(_13236_) );
	NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(_13235_), .B(_13236_), .C(_13234_), .Y(_13237_) );
	OAI22X1 OAI22X1_825 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_30_), .B(_13497_), .C(_13674_), .D(csr_gpr_iu_rs1_31_), .Y(_13238_) );
	INVX1 INVX1_2072 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .Y(_13239_) );
	OAI21X1 OAI21X1_5361 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_30_), .B(_12015_), .C(_13239_), .Y(_13240_) );
	NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_13238_), .B(_13240_), .Y(_13241_) );
	INVX1 INVX1_2073 ( .gnd(gnd), .vdd(vdd), .A(_13241_), .Y(_13242_) );
	XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_29_), .B(csr_gpr_iu_rs1_29_), .Y(_13243_) );
	XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(csr_gpr_iu_rs1_28_), .Y(_13244_) );
	NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_13244_), .B(_13243_), .Y(_13245_) );
	NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_13245_), .B(_13242_), .Y(_13246_) );
	OAI22X1 OAI22X1_826 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_26_), .B(_11887_), .C(_13508_), .D(csr_gpr_iu_rs1_27_), .Y(_13247_) );
	NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_27_), .B(_13508_), .Y(_13248_) );
	OAI21X1 OAI21X1_5362 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_26_), .B(_11884_), .C(_13248_), .Y(_13249_) );
	NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_13247_), .B(_13249_), .Y(_13250_) );
	NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_13250_), .B(_13246_), .Y(_13251_) );
	NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_13237_), .B(_13251_), .Y(_13252_) );
	INVX1 INVX1_2074 ( .gnd(gnd), .vdd(vdd), .A(_13252_), .Y(_13253_) );
	OAI22X1 OAI22X1_827 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_22_), .B(_13533_), .C(_13526_), .D(csr_gpr_iu_rs1_23_), .Y(_13254_) );
	NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_23_), .B(_13526_), .Y(_13255_) );
	OAI21X1 OAI21X1_5363 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_22_), .B(_11757_), .C(_13255_), .Y(_13256_) );
	NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .B(_13256_), .Y(_13257_) );
	INVX1 INVX1_2075 ( .gnd(gnd), .vdd(vdd), .A(_13257_), .Y(_13258_) );
	XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_21_), .B(csr_gpr_iu_rs1_21_), .Y(_13259_) );
	NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(csr_gpr_iu_rs1_20_), .Y(_13260_) );
	NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_11696_), .Y(_13261_) );
	OAI21X1 OAI21X1_5364 ( .gnd(gnd), .vdd(vdd), .A(_13260_), .B(_13261_), .C(_13259_), .Y(_13262_) );
	NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_13262_), .B(_13258_), .Y(_13263_) );
	OAI22X1 OAI22X1_828 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_18_), .B(_13550_), .C(_13545_), .D(csr_gpr_iu_rs1_19_), .Y(_13264_) );
	INVX1 INVX1_2076 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_18_), .Y(_13265_) );
	NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_19_), .B(_13545_), .Y(_13266_) );
	OAI21X1 OAI21X1_5365 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_18_), .B(_13265_), .C(_13266_), .Y(_13267_) );
	NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13267_), .Y(_13268_) );
	NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_11578_), .Y(_13269_) );
	NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(csr_gpr_iu_rs1_16_), .Y(_13270_) );
	NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_11604_), .Y(_13271_) );
	INVX1 INVX1_2077 ( .gnd(gnd), .vdd(vdd), .A(_13271_), .Y(_13272_) );
	NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_17_), .B(_11604_), .Y(_13273_) );
	NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_13273_), .B(_13272_), .Y(_13274_) );
	AOI21X1 AOI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_13269_), .B(_13270_), .C(_13274_), .Y(_13275_) );
	NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(_13268_), .B(_13275_), .C(_13263_), .Y(_13276_) );
	NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_13276_), .B(_13253_), .Y(_13277_) );
	OAI22X1 OAI22X1_829 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_14_), .B(_11499_), .C(_13570_), .D(csr_gpr_iu_rs1_15_), .Y(_13278_) );
	OAI22X1 OAI22X1_830 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_11540_), .C(csr_gpr_iu_rs2_14_), .D(_11504_), .Y(_13279_) );
	NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_13278_), .B(_13279_), .Y(_13280_) );
	INVX1 INVX1_2078 ( .gnd(gnd), .vdd(vdd), .A(_13280_), .Y(_13281_) );
	NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_13_), .B(_11469_), .Y(_13282_) );
	NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .B(_13577_), .Y(_13283_) );
	NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_13282_), .B(_13283_), .Y(_13284_) );
	NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .B(_13564_), .Y(_13285_) );
	NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_12_), .B(_11435_), .Y(_13286_) );
	NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(_13285_), .B(_13286_), .C(_13284_), .Y(_13287_) );
	NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_13281_), .B(_13287_), .Y(_13288_) );
	NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_8_), .B(_13980_), .Y(_13289_) );
	OAI21X1 OAI21X1_5366 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .B(_11322_), .C(_13289_), .Y(_13290_) );
	NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .B(_11322_), .Y(_13291_) );
	OAI21X1 OAI21X1_5367 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_8_), .B(_13980_), .C(_13291_), .Y(_13292_) );
	NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_13290_), .B(_13292_), .Y(_13293_) );
	OAI22X1 OAI22X1_831 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .B(_11351_), .C(_13587_), .D(csr_gpr_iu_rs1_11_), .Y(_13294_) );
	OAI22X1 OAI22X1_832 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_11390_), .C(csr_gpr_iu_rs2_10_), .D(_11356_), .Y(_13295_) );
	NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .B(_13295_), .Y(_13296_) );
	NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(_13293_), .B(_13296_), .C(_13288_), .Y(_13297_) );
	NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .B(_13885_), .Y(_13298_) );
	NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_7_), .B(_13640_), .Y(_13299_) );
	NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_7_), .B(_13927_), .Y(_13300_) );
	NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_13299_), .B(_13300_), .Y(_13301_) );
	OAI21X1 OAI21X1_5368 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_6_), .B(_13905_), .C(_13301_), .Y(_13302_) );
	OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_13302_), .B(_13298_), .Y(_13303_) );
	NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_5_), .B(_13854_), .Y(_13304_) );
	NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .B(_13612_), .Y(_13305_) );
	NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(_13305_), .Y(_13306_) );
	NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_4_), .B(csr_gpr_iu_rs1_4_), .Y(_13307_) );
	NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_13451_), .B(_13810_), .Y(_13308_) );
	OAI21X1 OAI21X1_5369 ( .gnd(gnd), .vdd(vdd), .A(_13307_), .B(_13308_), .C(_13306_), .Y(_13309_) );
	NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_13309_), .B(_13303_), .Y(_13310_) );
	NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .B(_13435_), .Y(_13311_) );
	NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_2_), .B(_13758_), .Y(_13312_) );
	NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .B(_13622_), .Y(_13313_) );
	NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .B(_13622_), .Y(_13314_) );
	INVX1 INVX1_2079 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .Y(_13315_) );
	NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_13313_), .B(_13315_), .Y(_13316_) );
	OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_13316_), .B(_13312_), .Y(_13317_) );
	NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_13311_), .B(_13317_), .Y(_13318_) );
	NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_1_), .B(_13705_), .Y(_13319_) );
	NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_1_), .B(_13630_), .Y(_13320_) );
	NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_13319_), .B(_13320_), .Y(_13321_) );
	OAI21X1 OAI21X1_5370 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_13455_), .C(_13321_), .Y(_13322_) );
	AOI21X1 AOI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(_13455_), .C(_13322_), .Y(_13323_) );
	NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(_13318_), .B(_13323_), .C(_13310_), .Y(_13324_) );
	NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_13297_), .B(_13324_), .Y(_13325_) );
	NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_13325_), .B(_13277_), .Y(_13326_) );
	AOI21X1 AOI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_13311_), .B(_13313_), .C(_13314_), .Y(_13327_) );
	OAI21X1 OAI21X1_5371 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(csr_gpr_iu_rs1_1_), .C(_13322_), .Y(_13328_) );
	NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_13318_), .B(_13328_), .Y(_13329_) );
	NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_13327_), .B(_13329_), .Y(_13330_) );
	NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_4_), .B(_13451_), .Y(_13331_) );
	AOI21X1 AOI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_13306_), .B(_13331_), .C(_13305_), .Y(_13332_) );
	AOI21X1 AOI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_13301_), .B(_13298_), .C(_13299_), .Y(_13333_) );
	OAI21X1 OAI21X1_5372 ( .gnd(gnd), .vdd(vdd), .A(_13332_), .B(_13303_), .C(_13333_), .Y(_13334_) );
	AOI21X1 AOI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_13330_), .B(_13310_), .C(_13334_), .Y(_13335_) );
	NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_9_), .B(_11322_), .Y(_13336_) );
	OAI21X1 OAI21X1_5373 ( .gnd(gnd), .vdd(vdd), .A(_13289_), .B(_13336_), .C(_13291_), .Y(_13337_) );
	NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_13337_), .B(_13296_), .Y(_13338_) );
	OAI21X1 OAI21X1_5374 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_11_), .B(_11390_), .C(_13294_), .Y(_13339_) );
	NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13338_), .Y(_13340_) );
	NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_13286_), .B(_13282_), .Y(_13341_) );
	OAI21X1 OAI21X1_5375 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .B(_13341_), .C(_13280_), .Y(_13342_) );
	OAI21X1 OAI21X1_5376 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_15_), .B(_11540_), .C(_13278_), .Y(_13343_) );
	NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_13343_), .B(_13342_), .Y(_13344_) );
	AOI21X1 AOI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_13288_), .B(_13340_), .C(_13344_), .Y(_13345_) );
	OAI21X1 OAI21X1_5377 ( .gnd(gnd), .vdd(vdd), .A(_13297_), .B(_13335_), .C(_13345_), .Y(_13346_) );
	NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_13346_), .Y(_13347_) );
	INVX1 INVX1_2080 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .Y(_13348_) );
	NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_16_), .B(_11578_), .Y(_13349_) );
	OAI21X1 OAI21X1_5378 ( .gnd(gnd), .vdd(vdd), .A(_13349_), .B(_13271_), .C(_13273_), .Y(_13350_) );
	AOI22X1 AOI22X1_679 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13266_), .C(_13350_), .D(_13268_), .Y(_13351_) );
	NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_20_), .B(_11696_), .C(_13259_), .Y(_13352_) );
	OAI21X1 OAI21X1_5379 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(csr_gpr_iu_rs1_21_), .C(_13352_), .Y(_13353_) );
	AOI22X1 AOI22X1_680 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .B(_13255_), .C(_13257_), .D(_13353_), .Y(_13354_) );
	OAI21X1 OAI21X1_5380 ( .gnd(gnd), .vdd(vdd), .A(_13351_), .B(_13348_), .C(_13354_), .Y(_13355_) );
	INVX1 INVX1_2081 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .Y(_13356_) );
	NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_28_), .B(_11951_), .C(_13243_), .Y(_13357_) );
	OAI21X1 OAI21X1_5381 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(csr_gpr_iu_rs1_29_), .C(_13357_), .Y(_13358_) );
	AOI22X1 AOI22X1_681 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13238_), .C(_13358_), .D(_13241_), .Y(_13359_) );
	INVX1 INVX1_2082 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .Y(_13360_) );
	OAI21X1 OAI21X1_5382 ( .gnd(gnd), .vdd(vdd), .A(_13236_), .B(_13232_), .C(_13360_), .Y(_13361_) );
	AOI22X1 AOI22X1_682 ( .gnd(gnd), .vdd(vdd), .A(_13247_), .B(_13248_), .C(_13361_), .D(_13250_), .Y(_13362_) );
	OAI21X1 OAI21X1_5383 ( .gnd(gnd), .vdd(vdd), .A(_13362_), .B(_13356_), .C(_13359_), .Y(_13363_) );
	AOI21X1 AOI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_13252_), .B(_13355_), .C(_13363_), .Y(_13364_) );
	NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_13364_), .B(_13347_), .Y(_13365_) );
	AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_13365_), .B(_13326_), .Y(_13366_) );
	NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(_13366_), .Y(_13367_) );
	OAI21X1 OAI21X1_5384 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_31_), .B(_13674_), .C(blt), .Y(_13368_) );
	INVX1 INVX1_2083 ( .gnd(gnd), .vdd(vdd), .A(bgeu), .Y(_13369_) );
	MUX2X1 MUX2X1_200 ( .gnd(gnd), .vdd(vdd), .A(bne), .B(beq), .S(_13326_), .Y(_13370_) );
	OAI21X1 OAI21X1_5385 ( .gnd(gnd), .vdd(vdd), .A(_13369_), .B(_13365_), .C(_13370_), .Y(_13371_) );
	NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_12337__bF_buf0), .B(_13371_), .Y(_13372_) );
	OAI21X1 OAI21X1_5386 ( .gnd(gnd), .vdd(vdd), .A(bge), .B(bltu), .C(_13366_), .Y(_13373_) );
	AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_13372_), .B(_13373_), .Y(_13374_) );
	OAI21X1 OAI21X1_5387 ( .gnd(gnd), .vdd(vdd), .A(_13367_), .B(_13368_), .C(_13374_), .Y(exu_alu_pc_jmp) );
	NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_0_), .B(csr_gpr_iu_rs2_1_), .Y(_13375_) );
	NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13451_), .C(_13375_), .Y(_13376_) );
	NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs2_3_), .B(_13376_), .Y(_13377_) );
	NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_20_bF_buf2), .B(biu_ins_21_bF_buf2), .Y(_13378_) );
	NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_22_bF_buf0), .B(biu_ins_23_), .Y(_13379_) );
	AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13450_), .Y(_13380_) );
	NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_13378_), .B(_13380_), .Y(_13381_) );
	NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_0_), .B(_13432_), .Y(_13382_) );
	NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_shift_counter_1_), .B(_13382_), .Y(_13383_) );
	AOI21X1 AOI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_13383_), .B(_13390_), .C(_13417_), .Y(_13384_) );
	OAI21X1 OAI21X1_5388 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .B(_13381_), .C(_13384_), .Y(_13385_) );
	AOI21X1 AOI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .B(_13377_), .C(_13385_), .Y(_13386_) );
	NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_13397__bF_buf1), .B(_13386_), .Y(csr_gpr_iu_rdy_exu) );
	DFFPOSX1 DFFPOSX1_1911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_11292__0_), .Q(data_rd_0_) );
	DFFPOSX1 DFFPOSX1_1912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_11292__1_), .Q(data_rd_1_) );
	DFFPOSX1 DFFPOSX1_1913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_11292__2_), .Q(data_rd_2_) );
	DFFPOSX1 DFFPOSX1_1914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_11292__3_), .Q(data_rd_3_) );
	DFFPOSX1 DFFPOSX1_1915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_11292__4_), .Q(data_rd_4_) );
	DFFPOSX1 DFFPOSX1_1916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_11292__5_), .Q(data_rd_5_) );
	DFFPOSX1 DFFPOSX1_1917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_11292__6_), .Q(data_rd_6_) );
	DFFPOSX1 DFFPOSX1_1918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_11292__7_), .Q(data_rd_7_) );
	DFFPOSX1 DFFPOSX1_1919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_11292__8_), .Q(data_rd_8_) );
	DFFPOSX1 DFFPOSX1_1920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_11292__9_), .Q(data_rd_9_) );
	DFFPOSX1 DFFPOSX1_1921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_11292__10_), .Q(data_rd_10_) );
	DFFPOSX1 DFFPOSX1_1922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_11292__11_), .Q(data_rd_11_) );
	DFFPOSX1 DFFPOSX1_1923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_11292__12_), .Q(data_rd_12_) );
	DFFPOSX1 DFFPOSX1_1924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_11292__13_), .Q(data_rd_13_) );
	DFFPOSX1 DFFPOSX1_1925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_11292__14_), .Q(data_rd_14_) );
	DFFPOSX1 DFFPOSX1_1926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_11292__15_), .Q(data_rd_15_) );
	DFFPOSX1 DFFPOSX1_1927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_11292__16_), .Q(data_rd_16_) );
	DFFPOSX1 DFFPOSX1_1928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_11292__17_), .Q(data_rd_17_) );
	DFFPOSX1 DFFPOSX1_1929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_11292__18_), .Q(data_rd_18_) );
	DFFPOSX1 DFFPOSX1_1930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_11292__19_), .Q(data_rd_19_) );
	DFFPOSX1 DFFPOSX1_1931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_11292__20_), .Q(data_rd_20_) );
	DFFPOSX1 DFFPOSX1_1932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_11292__21_), .Q(data_rd_21_) );
	DFFPOSX1 DFFPOSX1_1933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_11292__22_), .Q(data_rd_22_) );
	DFFPOSX1 DFFPOSX1_1934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_11292__23_), .Q(data_rd_23_) );
	DFFPOSX1 DFFPOSX1_1935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_11292__24_), .Q(data_rd_24_) );
	DFFPOSX1 DFFPOSX1_1936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_11292__25_), .Q(data_rd_25_) );
	DFFPOSX1 DFFPOSX1_1937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_11292__26_), .Q(data_rd_26_) );
	DFFPOSX1 DFFPOSX1_1938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_11292__27_), .Q(data_rd_27_) );
	DFFPOSX1 DFFPOSX1_1939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_11292__28_), .Q(data_rd_28_) );
	DFFPOSX1 DFFPOSX1_1940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_11292__29_), .Q(data_rd_29_) );
	DFFPOSX1 DFFPOSX1_1941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_11292__30_), .Q(data_rd_30_) );
	DFFPOSX1 DFFPOSX1_1942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_11292__31_), .Q(data_rd_31_) );
	DFFPOSX1 DFFPOSX1_1943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_11293__0_), .Q(biu_biu_data_in_0_) );
	DFFPOSX1 DFFPOSX1_1944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_11293__1_), .Q(biu_biu_data_in_1_) );
	DFFPOSX1 DFFPOSX1_1945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_11293__2_), .Q(biu_biu_data_in_2_) );
	DFFPOSX1 DFFPOSX1_1946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_11293__3_), .Q(biu_biu_data_in_3_) );
	DFFPOSX1 DFFPOSX1_1947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_11293__4_), .Q(biu_biu_data_in_4_) );
	DFFPOSX1 DFFPOSX1_1948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_11293__5_), .Q(biu_biu_data_in_5_) );
	DFFPOSX1 DFFPOSX1_1949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_11293__6_), .Q(biu_biu_data_in_6_) );
	DFFPOSX1 DFFPOSX1_1950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_11293__7_), .Q(biu_biu_data_in_7_) );
	DFFPOSX1 DFFPOSX1_1951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_11293__8_), .Q(biu_biu_data_in_8_) );
	DFFPOSX1 DFFPOSX1_1952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_11293__9_), .Q(biu_biu_data_in_9_) );
	DFFPOSX1 DFFPOSX1_1953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_11293__10_), .Q(biu_biu_data_in_10_) );
	DFFPOSX1 DFFPOSX1_1954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_11293__11_), .Q(biu_biu_data_in_11_) );
	DFFPOSX1 DFFPOSX1_1955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_11293__12_), .Q(biu_biu_data_in_12_) );
	DFFPOSX1 DFFPOSX1_1956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_11293__13_), .Q(biu_biu_data_in_13_) );
	DFFPOSX1 DFFPOSX1_1957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_11293__14_), .Q(biu_biu_data_in_14_) );
	DFFPOSX1 DFFPOSX1_1958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_11293__15_), .Q(biu_biu_data_in_15_) );
	DFFPOSX1 DFFPOSX1_1959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_11293__16_), .Q(biu_biu_data_in_16_) );
	DFFPOSX1 DFFPOSX1_1960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_11293__17_), .Q(biu_biu_data_in_17_) );
	DFFPOSX1 DFFPOSX1_1961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_11293__18_), .Q(biu_biu_data_in_18_) );
	DFFPOSX1 DFFPOSX1_1962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_11293__19_), .Q(biu_biu_data_in_19_) );
	DFFPOSX1 DFFPOSX1_1963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_11293__20_), .Q(biu_biu_data_in_20_) );
	DFFPOSX1 DFFPOSX1_1964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_11293__21_), .Q(biu_biu_data_in_21_) );
	DFFPOSX1 DFFPOSX1_1965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_11293__22_), .Q(biu_biu_data_in_22_) );
	DFFPOSX1 DFFPOSX1_1966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_11293__23_), .Q(biu_biu_data_in_23_) );
	DFFPOSX1 DFFPOSX1_1967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_11293__24_), .Q(biu_biu_data_in_24_) );
	DFFPOSX1 DFFPOSX1_1968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_11293__25_), .Q(biu_biu_data_in_25_) );
	DFFPOSX1 DFFPOSX1_1969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_11293__26_), .Q(biu_biu_data_in_26_) );
	DFFPOSX1 DFFPOSX1_1970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_11293__27_), .Q(biu_biu_data_in_27_) );
	DFFPOSX1 DFFPOSX1_1971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_11293__28_), .Q(biu_biu_data_in_28_) );
	DFFPOSX1 DFFPOSX1_1972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_11293__29_), .Q(biu_biu_data_in_29_) );
	DFFPOSX1 DFFPOSX1_1973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_11293__30_), .Q(biu_biu_data_in_30_) );
	DFFPOSX1 DFFPOSX1_1974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_11293__31_), .Q(biu_biu_data_in_31_) );
	DFFPOSX1 DFFPOSX1_1975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_11294__0_), .Q(exu_alu_shift_counter_0_) );
	DFFPOSX1 DFFPOSX1_1976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_11294__1_), .Q(exu_alu_shift_counter_1_) );
	DFFPOSX1 DFFPOSX1_1977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_11294__2_), .Q(exu_alu_shift_counter_2_) );
	DFFPOSX1 DFFPOSX1_1978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_11294__3_), .Q(exu_alu_shift_counter_3_) );
	DFFPOSX1 DFFPOSX1_1979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_11294__4_), .Q(exu_alu_shift_counter_4_) );
	OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_2_), .B(biu_exce_chk_statu_cpu_1_), .Y(_14321_) );
	INVX1 INVX1_2084 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_3_), .Y(_14322_) );
	NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_statu_cpu_0_), .B(csr_gpr_iu_rdy_exu), .C(_14322_), .Y(_14323_) );
	NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf3), .B(_14323__bF_buf3), .Y(_14324_) );
	INVX2 INVX2_189 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .Y(_14325_) );
	NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14325_), .Y(_14326_) );
	MUX2X1 MUX2X1_201 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_0_), .B(csr_gpr_iu_rs1_0_), .S(_14326_), .Y(_14327_) );
	INVX8 INVX8_105 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf49), .Y(_14328_) );
	OAI21X1 OAI21X1_5389 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_0_), .B(_14324__bF_buf8), .C(_14328__bF_buf5), .Y(_14329_) );
	AOI21X1 AOI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_14324__bF_buf7), .B(_14327_), .C(_14329_), .Y(_13986__0_) );
	INVX1 INVX1_2085 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_1_), .Y(_14330_) );
	NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_ins_dec_jal_bF_buf3), .Y(_14331_) );
	INVX4 INVX4_60 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf3), .Y(_14332_) );
	INVX2 INVX2_190 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .Y(_14333_) );
	NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(_14333_), .Y(_14334_) );
	AOI22X1 AOI22X1_683 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_ins_12_), .C(csr_gpr_iu_imm12_0_), .D(_14334__bF_buf4), .Y(_14335_) );
	OAI21X1 OAI21X1_5390 ( .gnd(gnd), .vdd(vdd), .A(_14330_), .B(_14332_), .C(_14335_), .Y(_14336_) );
	NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(bne), .B(beq), .Y(_14337_) );
	NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(bltu), .B(blt), .Y(_14338_) );
	NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(bgeu), .B(bge), .Y(_14339_) );
	NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(_14337_), .B(_14338_), .C(_14339_), .Y(_14340_) );
	NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14340_), .Y(_14341_) );
	NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_0_), .B(_14331__bF_buf2), .Y(_14342_) );
	AOI22X1 AOI22X1_684 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_pc_1_), .C(csr_gpr_iu_rs1_1_), .D(_14334__bF_buf3), .Y(_14343_) );
	OAI21X1 OAI21X1_5391 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .B(_14341_), .C(_14343_), .Y(_14344_) );
	XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_14344_), .B(_14336_), .Y(_14345_) );
	OAI21X1 OAI21X1_5392 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_1_), .B(_14324__bF_buf6), .C(_14328__bF_buf4), .Y(_14346_) );
	AOI21X1 AOI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_14345_), .B(_14324__bF_buf5), .C(_14346_), .Y(_13986__1_) );
	NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_14336_), .B(_14344_), .Y(_14347_) );
	AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf1), .B(biu_pc_2_), .Y(_14348_) );
	INVX1 INVX1_2086 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_1_), .Y(_14349_) );
	NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_ins_13_), .Y(_14350_) );
	OAI21X1 OAI21X1_5393 ( .gnd(gnd), .vdd(vdd), .A(_14349_), .B(_14326_), .C(_14350_), .Y(_14351_) );
	NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_14348_), .B(_14351_), .Y(_14352_) );
	NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_pc_2_), .Y(_14353_) );
	INVX1 INVX1_2087 ( .gnd(gnd), .vdd(vdd), .A(_14353_), .Y(_14354_) );
	NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_imm12_1_), .Y(_14355_) );
	NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14355_), .C(_14340_), .Y(_14356_) );
	INVX2 INVX2_191 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .Y(_14357_) );
	AOI21X1 AOI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(csr_gpr_iu_ins_dec_jalr), .C(csr_gpr_iu_ins_dec_jal_bF_buf5), .Y(_14358_) );
	AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_14356_), .B(_14358_), .Y(_14359_) );
	OAI21X1 OAI21X1_5394 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .B(_14359_), .C(_14352_), .Y(_14360_) );
	INVX1 INVX1_2088 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .Y(_14361_) );
	NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14356_), .Y(_14362_) );
	NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(_14353_), .B(_14362_), .C(_14361_), .Y(_14363_) );
	AOI21X1 AOI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_14360_), .B(_14363_), .C(_14347_), .Y(_14364_) );
	INVX1 INVX1_2089 ( .gnd(gnd), .vdd(vdd), .A(_14364_), .Y(_14365_) );
	NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(_14347_), .B(_14363_), .C(_14360_), .Y(_14366_) );
	NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_14366_), .B(_14365_), .Y(_14367_) );
	OAI21X1 OAI21X1_5395 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_2_), .B(_14324__bF_buf4), .C(_14328__bF_buf3), .Y(_14368_) );
	AOI21X1 AOI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_14367_), .B(_14324__bF_buf3), .C(_14368_), .Y(_13986__2_) );
	NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .B(_14359_), .Y(_14369_) );
	OAI21X1 OAI21X1_5396 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .B(_14369_), .C(_14365_), .Y(_14370_) );
	INVX1 INVX1_2090 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .Y(_14371_) );
	NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(biu_ins_14_), .Y(_14372_) );
	OAI21X1 OAI21X1_5397 ( .gnd(gnd), .vdd(vdd), .A(_14371_), .B(_14326_), .C(_14372_), .Y(_14373_) );
	AOI21X1 AOI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_3_), .B(_14331__bF_buf0), .C(_14373_), .Y(_14374_) );
	AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_14340_), .B(exu_alu_pc_jmp), .Y(_14375_) );
	NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_2_), .B(_14331__bF_buf3), .C(_14375_), .Y(_14376_) );
	AOI22X1 AOI22X1_685 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(biu_pc_3_), .C(csr_gpr_iu_rs1_3_), .D(_14334__bF_buf2), .Y(_14377_) );
	AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_14376_), .B(_14377_), .Y(_14378_) );
	NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_14374_), .B(_14378_), .Y(_14379_) );
	OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_14378_), .B(_14374_), .Y(_14380_) );
	NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_14379_), .B(_14380_), .Y(_14381_) );
	XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_14370_), .B(_14381_), .Y(_14382_) );
	OAI21X1 OAI21X1_5398 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_3_), .B(_14324__bF_buf2), .C(_14328__bF_buf2), .Y(_14383_) );
	AOI21X1 AOI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_14382_), .B(_14324__bF_buf1), .C(_14383_), .Y(_13986__3_) );
	AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf2), .B(biu_pc_4_), .Y(_14384_) );
	INVX1 INVX1_2091 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_3_), .Y(_14385_) );
	NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_ins_15_bF_buf3), .Y(_14386_) );
	OAI21X1 OAI21X1_5399 ( .gnd(gnd), .vdd(vdd), .A(_14385_), .B(_14326_), .C(_14386_), .Y(_14387_) );
	NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_14384_), .B(_14387_), .Y(_14388_) );
	NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_14385_), .B(_14332_), .Y(_14389_) );
	NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_14389_), .B(_14375_), .Y(_14390_) );
	AOI22X1 AOI22X1_686 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_pc_4_), .C(csr_gpr_iu_rs1_4_), .D(_14334__bF_buf1), .Y(_14391_) );
	NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(_14388_), .B(_14391_), .C(_14390_), .Y(_14392_) );
	INVX1 INVX1_2092 ( .gnd(gnd), .vdd(vdd), .A(_14389_), .Y(_14393_) );
	OAI21X1 OAI21X1_5400 ( .gnd(gnd), .vdd(vdd), .A(_14341_), .B(_14393_), .C(_14391_), .Y(_14394_) );
	OAI21X1 OAI21X1_5401 ( .gnd(gnd), .vdd(vdd), .A(_14384_), .B(_14387_), .C(_14394_), .Y(_14395_) );
	AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .B(_14392_), .Y(_14396_) );
	INVX1 INVX1_2093 ( .gnd(gnd), .vdd(vdd), .A(_14396_), .Y(_14397_) );
	OAI22X1 OAI22X1_833 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .B(_14369_), .C(_14374_), .D(_14378_), .Y(_14398_) );
	OAI21X1 OAI21X1_5402 ( .gnd(gnd), .vdd(vdd), .A(_14398_), .B(_14364_), .C(_14379_), .Y(_14399_) );
	XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_14399_), .B(_14397_), .Y(_14400_) );
	OAI21X1 OAI21X1_5403 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_4_), .B(_14324__bF_buf0), .C(_14328__bF_buf1), .Y(_14401_) );
	AOI21X1 AOI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_14400_), .B(_14324__bF_buf8), .C(_14401_), .Y(_13986__4_) );
	OAI21X1 OAI21X1_5404 ( .gnd(gnd), .vdd(vdd), .A(_14397_), .B(_14399_), .C(_14395_), .Y(_14402_) );
	AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf1), .B(biu_pc_5_), .Y(_14403_) );
	INVX1 INVX1_2094 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_4_), .Y(_14404_) );
	NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_ins_16_), .Y(_14405_) );
	OAI21X1 OAI21X1_5405 ( .gnd(gnd), .vdd(vdd), .A(_14404_), .B(_14326_), .C(_14405_), .Y(_14406_) );
	NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_14403_), .B(_14406_), .Y(_14407_) );
	NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_imm12_4_), .B(_14331__bF_buf0), .Y(_14408_) );
	INVX1 INVX1_2095 ( .gnd(gnd), .vdd(vdd), .A(_14408_), .Y(_14409_) );
	NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14340_), .C(_14409_), .Y(_14410_) );
	AOI22X1 AOI22X1_687 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_pc_5_), .C(csr_gpr_iu_rs1_5_), .D(_14334__bF_buf0), .Y(_14411_) );
	NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(_14411_), .B(_14410_), .C(_14407_), .Y(_14412_) );
	OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_14406_), .B(_14403_), .Y(_14413_) );
	OAI21X1 OAI21X1_5406 ( .gnd(gnd), .vdd(vdd), .A(_14408_), .B(_14341_), .C(_14411_), .Y(_14414_) );
	NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_14413_), .B(_14414_), .Y(_14415_) );
	NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_14412_), .B(_14415_), .Y(_14416_) );
	INVX2 INVX2_192 ( .gnd(gnd), .vdd(vdd), .A(_14416_), .Y(_14417_) );
	XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_14402_), .B(_14417_), .Y(_14418_) );
	OAI21X1 OAI21X1_5407 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_5_), .B(_14324__bF_buf7), .C(_14328__bF_buf0), .Y(_14419_) );
	AOI21X1 AOI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_14418_), .B(_14324__bF_buf6), .C(_14419_), .Y(_13986__5_) );
	NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_14417_), .B(_14396_), .Y(_14420_) );
	OAI21X1 OAI21X1_5408 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .B(_14416_), .C(_14415_), .Y(_14421_) );
	INVX1 INVX1_2096 ( .gnd(gnd), .vdd(vdd), .A(_14421_), .Y(_14422_) );
	OAI21X1 OAI21X1_5409 ( .gnd(gnd), .vdd(vdd), .A(_14420_), .B(_14399_), .C(_14422_), .Y(_14423_) );
	AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf3), .B(biu_pc_6_), .Y(_14424_) );
	INVX1 INVX1_2097 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf3), .Y(_14425_) );
	NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_ins_17_), .Y(_14426_) );
	OAI21X1 OAI21X1_5410 ( .gnd(gnd), .vdd(vdd), .A(_14425_), .B(_14326_), .C(_14426_), .Y(_14427_) );
	NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_14424_), .B(_14427_), .Y(_14428_) );
	NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_25_bF_buf2), .B(_14331__bF_buf2), .Y(_14429_) );
	AOI22X1 AOI22X1_688 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(biu_pc_6_), .C(csr_gpr_iu_rs1_6_), .D(_14334__bF_buf4), .Y(_14430_) );
	OAI21X1 OAI21X1_5411 ( .gnd(gnd), .vdd(vdd), .A(_14429_), .B(_14341_), .C(_14430_), .Y(_14431_) );
	NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_14428_), .B(_14431_), .Y(_14432_) );
	OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_14431_), .B(_14428_), .Y(_14433_) );
	NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_14432_), .B(_14433_), .Y(_14434_) );
	XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14434_), .Y(_14435_) );
	OAI21X1 OAI21X1_5412 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_6_), .B(_14324__bF_buf5), .C(_14328__bF_buf5), .Y(_14436_) );
	AOI21X1 AOI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_14435_), .B(_14324__bF_buf4), .C(_14436_), .Y(_13986__6_) );
	OAI21X1 OAI21X1_5413 ( .gnd(gnd), .vdd(vdd), .A(_14424_), .B(_14427_), .C(_14431_), .Y(_14437_) );
	INVX1 INVX1_2098 ( .gnd(gnd), .vdd(vdd), .A(_14437_), .Y(_14438_) );
	AOI21X1 AOI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14434_), .C(_14438_), .Y(_14439_) );
	AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf1), .B(biu_pc_7_), .Y(_14440_) );
	INVX1 INVX1_2099 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf1), .Y(_14441_) );
	NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(biu_ins_18_), .Y(_14442_) );
	OAI21X1 OAI21X1_5414 ( .gnd(gnd), .vdd(vdd), .A(_14441_), .B(_14326_), .C(_14442_), .Y(_14443_) );
	NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_14440_), .B(_14443_), .Y(_14444_) );
	NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_26_bF_buf0), .B(_14331__bF_buf0), .Y(_14445_) );
	INVX1 INVX1_2100 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .Y(_14446_) );
	NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14340_), .C(_14446_), .Y(_14447_) );
	AOI22X1 AOI22X1_689 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(biu_pc_7_), .C(csr_gpr_iu_rs1_7_), .D(_14334__bF_buf3), .Y(_14448_) );
	NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(_14448_), .B(_14447_), .C(_14444_), .Y(_14449_) );
	OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_14443_), .B(_14440_), .Y(_14450_) );
	OAI21X1 OAI21X1_5415 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .B(_14341_), .C(_14448_), .Y(_14451_) );
	NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_14450_), .B(_14451_), .Y(_14452_) );
	NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_14449_), .B(_14452_), .Y(_14453_) );
	XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_14439_), .B(_14453_), .Y(_14454_) );
	OAI21X1 OAI21X1_5416 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_7_), .B(_14324__bF_buf3), .C(_14328__bF_buf4), .Y(_14455_) );
	AOI21X1 AOI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_14454_), .B(_14324__bF_buf2), .C(_14455_), .Y(_13986__7_) );
	AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf3), .B(biu_pc_8_), .Y(_14456_) );
	INVX1 INVX1_2101 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf0), .Y(_14457_) );
	NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_ins_19_), .Y(_14458_) );
	OAI21X1 OAI21X1_5417 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_14326_), .C(_14458_), .Y(_14459_) );
	NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_14456_), .B(_14459_), .Y(_14460_) );
	NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_27_bF_buf3), .B(_14331__bF_buf2), .Y(_14461_) );
	AOI22X1 AOI22X1_690 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_pc_8_), .C(csr_gpr_iu_rs1_8_), .D(_14334__bF_buf2), .Y(_14462_) );
	OAI21X1 OAI21X1_5418 ( .gnd(gnd), .vdd(vdd), .A(_14461_), .B(_14341_), .C(_14462_), .Y(_14463_) );
	NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_14460_), .B(_14463_), .Y(_14464_) );
	OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_14463_), .B(_14460_), .Y(_14465_) );
	NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_14464_), .B(_14465_), .Y(_14466_) );
	NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_14452_), .B(_14437_), .Y(_14467_) );
	AOI21X1 AOI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_14432_), .B(_14433_), .C(_14453_), .Y(_14468_) );
	AOI22X1 AOI22X1_691 ( .gnd(gnd), .vdd(vdd), .A(_14449_), .B(_14467_), .C(_14468_), .D(_14421_), .Y(_14469_) );
	NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(_14417_), .B(_14396_), .C(_14468_), .Y(_14470_) );
	OAI21X1 OAI21X1_5419 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14399_), .C(_14469_), .Y(_14471_) );
	XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_14471_), .B(_14466_), .Y(_14472_) );
	OAI21X1 OAI21X1_5420 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_8_), .B(_14324__bF_buf1), .C(_14328__bF_buf3), .Y(_14473_) );
	AOI21X1 AOI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_14472_), .B(_14324__bF_buf0), .C(_14473_), .Y(_13986__8_) );
	OAI21X1 OAI21X1_5421 ( .gnd(gnd), .vdd(vdd), .A(_14456_), .B(_14459_), .C(_14463_), .Y(_14474_) );
	INVX1 INVX1_2102 ( .gnd(gnd), .vdd(vdd), .A(_14474_), .Y(_14475_) );
	AOI21X1 AOI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_14471_), .B(_14466_), .C(_14475_), .Y(_14476_) );
	AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf1), .B(biu_pc_9_), .Y(_14477_) );
	INVX1 INVX1_2103 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf1), .Y(_14478_) );
	NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_ins_20_bF_buf1), .Y(_14479_) );
	OAI21X1 OAI21X1_5422 ( .gnd(gnd), .vdd(vdd), .A(_14478_), .B(_14326_), .C(_14479_), .Y(_14480_) );
	NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_14477_), .B(_14480_), .Y(_14481_) );
	NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_28_bF_buf0), .B(_14331__bF_buf0), .Y(_14482_) );
	INVX1 INVX1_2104 ( .gnd(gnd), .vdd(vdd), .A(_14482_), .Y(_14483_) );
	NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14340_), .C(_14483_), .Y(_14484_) );
	AOI22X1 AOI22X1_692 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_pc_9_), .C(csr_gpr_iu_rs1_9_), .D(_14334__bF_buf1), .Y(_14485_) );
	NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(_14485_), .B(_14484_), .C(_14481_), .Y(_14486_) );
	OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_14480_), .B(_14477_), .Y(_14487_) );
	OAI21X1 OAI21X1_5423 ( .gnd(gnd), .vdd(vdd), .A(_14482_), .B(_14341_), .C(_14485_), .Y(_14488_) );
	NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_14487_), .B(_14488_), .Y(_14489_) );
	NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_14486_), .B(_14489_), .Y(_14490_) );
	XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_14476_), .B(_14490_), .Y(_14491_) );
	OAI21X1 OAI21X1_5424 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_9_), .B(_14324__bF_buf8), .C(_14328__bF_buf2), .Y(_14492_) );
	AOI21X1 AOI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_14491_), .B(_14324__bF_buf7), .C(_14492_), .Y(_13986__9_) );
	INVX1 INVX1_2105 ( .gnd(gnd), .vdd(vdd), .A(_14486_), .Y(_14493_) );
	OAI21X1 OAI21X1_5425 ( .gnd(gnd), .vdd(vdd), .A(_14474_), .B(_14493_), .C(_14489_), .Y(_14494_) );
	INVX1 INVX1_2106 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .Y(_14495_) );
	AOI21X1 AOI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_14464_), .B(_14465_), .C(_14490_), .Y(_14496_) );
	NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14471_), .Y(_14497_) );
	NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_14495_), .B(_14497_), .Y(_14498_) );
	AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf3), .B(biu_pc_10_), .Y(_14499_) );
	INVX1 INVX1_2107 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_29_bF_buf2), .Y(_14500_) );
	NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_ins_21_bF_buf1), .Y(_14501_) );
	OAI21X1 OAI21X1_5426 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14326_), .C(_14501_), .Y(_14502_) );
	NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_14499_), .B(_14502_), .Y(_14503_) );
	NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_ins_dec_jal_bF_buf5), .C(_14500_), .Y(_14504_) );
	NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14504_), .C(_14340_), .Y(_14505_) );
	AOI22X1 AOI22X1_693 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(biu_pc_10_), .C(csr_gpr_iu_rs1_10_), .D(_14334__bF_buf0), .Y(_14506_) );
	NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(_14505_), .B(_14506_), .C(_14503_), .Y(_14507_) );
	NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_14506_), .B(_14505_), .Y(_14508_) );
	OAI21X1 OAI21X1_5427 ( .gnd(gnd), .vdd(vdd), .A(_14499_), .B(_14502_), .C(_14508_), .Y(_14509_) );
	NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_14507_), .B(_14509_), .Y(_14510_) );
	INVX1 INVX1_2108 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .Y(_14511_) );
	XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_14498_), .B(_14511_), .Y(_14512_) );
	OAI21X1 OAI21X1_5428 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_10_), .B(_14324__bF_buf6), .C(_14328__bF_buf1), .Y(_14513_) );
	AOI21X1 AOI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_14512_), .B(_14324__bF_buf5), .C(_14513_), .Y(_13986__10_) );
	NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .B(_14498_), .Y(_14514_) );
	NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_14509_), .B(_14514_), .Y(_14515_) );
	AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf2), .B(biu_pc_11_), .Y(_14516_) );
	INVX1 INVX1_2109 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_30_bF_buf0), .Y(_14517_) );
	NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(biu_ins_22_bF_buf3), .Y(_14518_) );
	OAI21X1 OAI21X1_5429 ( .gnd(gnd), .vdd(vdd), .A(_14517_), .B(_14326_), .C(_14518_), .Y(_14519_) );
	NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_14516_), .B(_14519_), .Y(_14520_) );
	AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_14331__bF_buf1), .B(biu_ins_30_bF_buf3), .Y(_14521_) );
	NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14340_), .C(_14521_), .Y(_14522_) );
	AOI22X1 AOI22X1_694 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_pc_11_), .C(csr_gpr_iu_rs1_11_), .D(_14334__bF_buf4), .Y(_14523_) );
	NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(_14522_), .B(_14523_), .C(_14520_), .Y(_14524_) );
	NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_14523_), .B(_14522_), .Y(_14525_) );
	OAI21X1 OAI21X1_5430 ( .gnd(gnd), .vdd(vdd), .A(_14516_), .B(_14519_), .C(_14525_), .Y(_14526_) );
	NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_14524_), .B(_14526_), .Y(_14527_) );
	XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_14515_), .B(_14527_), .Y(_14528_) );
	OAI21X1 OAI21X1_5431 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_11_), .B(_14324__bF_buf4), .C(_14328__bF_buf0), .Y(_14529_) );
	AOI21X1 AOI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_14528_), .B(_14324__bF_buf3), .C(_14529_), .Y(_13986__11_) );
	NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .B(_14527_), .Y(_14530_) );
	OAI21X1 OAI21X1_5432 ( .gnd(gnd), .vdd(vdd), .A(_14509_), .B(_14527_), .C(_14526_), .Y(_14531_) );
	AOI21X1 AOI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_14530_), .B(_14494_), .C(_14531_), .Y(_14532_) );
	NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14530_), .C(_14471_), .Y(_14533_) );
	NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_14532_), .B(_14533_), .Y(_14534_) );
	NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(_14331__bF_buf0), .C(_14375_), .Y(_14535_) );
	AOI22X1 AOI22X1_695 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_pc_12_), .C(csr_gpr_iu_rs1_12_), .D(_14334__bF_buf3), .Y(_14536_) );
	NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_12_), .B(_14333_), .Y(_14537_) );
	NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(biu_ins_31_bF_buf2), .Y(_14538_) );
	AOI21X1 AOI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_14537_), .B(_14538_), .C(csr_gpr_iu_ins_dec_jal_bF_buf0), .Y(_14539_) );
	AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_ins_23_), .Y(_14540_) );
	NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_14540_), .B(_14539_), .Y(_14541_) );
	NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(_14536_), .B(_14541_), .C(_14535_), .Y(_14542_) );
	INVX4 INVX4_61 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .Y(_14543_) );
	NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14543_), .Y(_14544_) );
	NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(exu_alu_pc_jmp), .B(_14544_), .C(_14340_), .Y(_14545_) );
	OAI21X1 OAI21X1_5433 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(_14545__bF_buf3), .C(_14536_), .Y(_14546_) );
	OAI21X1 OAI21X1_5434 ( .gnd(gnd), .vdd(vdd), .A(_14539_), .B(_14540_), .C(_14546_), .Y(_14547_) );
	AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_14542_), .B(_14547_), .Y(_14548_) );
	XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_14534_), .B(_14548_), .Y(_14549_) );
	OAI21X1 OAI21X1_5435 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_12_), .B(_14324__bF_buf2), .C(_14328__bF_buf5), .Y(_14550_) );
	AOI21X1 AOI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_14549_), .B(_14324__bF_buf1), .C(_14550_), .Y(_13986__12_) );
	INVX1 INVX1_2110 ( .gnd(gnd), .vdd(vdd), .A(_14534_), .Y(_14551_) );
	NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14542_), .Y(_14552_) );
	OAI21X1 OAI21X1_5436 ( .gnd(gnd), .vdd(vdd), .A(_14552_), .B(_14551_), .C(_14547_), .Y(_14553_) );
	AOI22X1 AOI22X1_696 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(biu_pc_13_), .C(csr_gpr_iu_rs1_13_), .D(_14334__bF_buf2), .Y(_14554_) );
	OAI21X1 OAI21X1_5437 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(_14545__bF_buf2), .C(_14554_), .Y(_14555_) );
	INVX1 INVX1_2111 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_24_), .Y(_14556_) );
	INVX1 INVX1_2112 ( .gnd(gnd), .vdd(vdd), .A(_14538_), .Y(_14557_) );
	NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(_14557_), .Y(_14558_) );
	NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_13_), .B(_14333_), .Y(_14559_) );
	AOI22X1 AOI22X1_697 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(_14556_), .C(_14559_), .D(_14558_), .Y(_14560_) );
	NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_14560_), .B(_14555_), .Y(_14561_) );
	AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_14555_), .B(_14560_), .Y(_14562_) );
	NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .B(_14562_), .Y(_14563_) );
	XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14553_), .B(_14563_), .Y(_14564_) );
	OAI21X1 OAI21X1_5438 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_13_), .B(_14324__bF_buf0), .C(_14328__bF_buf4), .Y(_14565_) );
	AOI21X1 AOI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_14564_), .B(_14324__bF_buf8), .C(_14565_), .Y(_13986__13_) );
	NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_14560_), .B(_14555_), .Y(_14566_) );
	OAI21X1 OAI21X1_5439 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14561_), .C(_14566_), .Y(_14567_) );
	XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_14555_), .B(_14560_), .Y(_14568_) );
	NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_14552_), .B(_14568_), .Y(_14569_) );
	AOI21X1 AOI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_14534_), .B(_14569_), .C(_14567_), .Y(_14570_) );
	AOI22X1 AOI22X1_698 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_pc_14_), .C(csr_gpr_iu_rs1_14_), .D(_14334__bF_buf1), .Y(_14571_) );
	OAI21X1 OAI21X1_5440 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(_14545__bF_buf1), .C(_14571_), .Y(_14572_) );
	NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_14_), .B(_14333_), .Y(_14573_) );
	NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_14573_), .B(_14558_), .Y(_14574_) );
	OAI21X1 OAI21X1_5441 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(biu_ins_25_bF_buf1), .C(_14574_), .Y(_14575_) );
	NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_14575_), .B(_14572_), .Y(_14576_) );
	OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_14572_), .B(_14575_), .Y(_14577_) );
	NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_14576_), .B(_14577_), .Y(_14578_) );
	INVX1 INVX1_2113 ( .gnd(gnd), .vdd(vdd), .A(_14578_), .Y(_14579_) );
	XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_14570_), .B(_14579_), .Y(_14580_) );
	OAI21X1 OAI21X1_5442 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_14_), .B(_14324__bF_buf7), .C(_14328__bF_buf3), .Y(_14581_) );
	AOI21X1 AOI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14324__bF_buf6), .C(_14581_), .Y(_13986__14_) );
	INVX1 INVX1_2114 ( .gnd(gnd), .vdd(vdd), .A(_14575_), .Y(_14582_) );
	NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_14572_), .B(_14582_), .Y(_14583_) );
	OAI21X1 OAI21X1_5443 ( .gnd(gnd), .vdd(vdd), .A(_14579_), .B(_14570_), .C(_14583_), .Y(_14584_) );
	AOI22X1 AOI22X1_699 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_pc_15_), .C(csr_gpr_iu_rs1_15_), .D(_14334__bF_buf0), .Y(_14585_) );
	NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_15_), .B(_14333_), .Y(_14586_) );
	AOI21X1 AOI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_14586_), .B(_14538_), .C(csr_gpr_iu_ins_dec_jal_bF_buf6), .Y(_14587_) );
	AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(biu_ins_26_bF_buf3), .Y(_14588_) );
	NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_14588_), .B(_14587_), .Y(_14589_) );
	NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(_14585_), .B(_14589_), .C(_14535_), .Y(_14590_) );
	OAI21X1 OAI21X1_5444 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(_14545__bF_buf0), .C(_14585_), .Y(_14591_) );
	OAI21X1 OAI21X1_5445 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .B(_14588_), .C(_14591_), .Y(_14592_) );
	AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_14590_), .B(_14592_), .Y(_14593_) );
	XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_14584_), .B(_14593_), .Y(_14594_) );
	OAI21X1 OAI21X1_5446 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_15_), .B(_14324__bF_buf5), .C(_14328__bF_buf2), .Y(_14595_) );
	AOI21X1 AOI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_14594_), .B(_14324__bF_buf4), .C(_14595_), .Y(_13986__15_) );
	NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_14530_), .B(_14496_), .Y(_14596_) );
	NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_14548_), .B(_14563_), .Y(_14597_) );
	NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_14593_), .B(_14578_), .Y(_14598_) );
	NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .B(_14598_), .C(_14596_), .Y(_14599_) );
	NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_14592_), .B(_14590_), .Y(_14600_) );
	AOI21X1 AOI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_14576_), .B(_14577_), .C(_14600_), .Y(_14601_) );
	NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14569_), .Y(_14602_) );
	OAI21X1 OAI21X1_5447 ( .gnd(gnd), .vdd(vdd), .A(_14583_), .B(_14600_), .C(_14592_), .Y(_14603_) );
	AOI21X1 AOI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14567_), .C(_14603_), .Y(_14604_) );
	OAI21X1 OAI21X1_5448 ( .gnd(gnd), .vdd(vdd), .A(_14532_), .B(_14602_), .C(_14604_), .Y(_14605_) );
	AOI21X1 AOI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_14471_), .B(_14599_), .C(_14605_), .Y(_14606_) );
	AOI22X1 AOI22X1_700 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(biu_pc_16_), .C(csr_gpr_iu_rs1_16_), .D(_14334__bF_buf4), .Y(_14607_) );
	OAI21X1 OAI21X1_5449 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(_14545__bF_buf3), .C(_14607_), .Y(_14608_) );
	INVX1 INVX1_2115 ( .gnd(gnd), .vdd(vdd), .A(_14608_), .Y(_14609_) );
	INVX1 INVX1_2116 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_16_), .Y(_14610_) );
	OAI21X1 OAI21X1_5450 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14610_), .C(_14558_), .Y(_14611_) );
	OAI21X1 OAI21X1_5451 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(biu_ins_27_bF_buf2), .C(_14611_), .Y(_14612_) );
	NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_14612_), .B(_14609_), .Y(_14613_) );
	OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_14609_), .B(_14612_), .Y(_14614_) );
	NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_14613_), .B(_14614_), .Y(_14615_) );
	XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_14606_), .B(_14615_), .Y(_14616_) );
	OAI21X1 OAI21X1_5452 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_16_), .B(_14324__bF_buf3), .C(_14328__bF_buf1), .Y(_14617_) );
	AOI21X1 AOI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_14616_), .B(_14324__bF_buf2), .C(_14617_), .Y(_13986__16_) );
	OAI21X1 OAI21X1_5453 ( .gnd(gnd), .vdd(vdd), .A(_14615_), .B(_14606_), .C(_14614_), .Y(_14618_) );
	AOI22X1 AOI22X1_701 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(biu_pc_17_), .C(csr_gpr_iu_rs1_17_), .D(_14334__bF_buf3), .Y(_14619_) );
	OAI21X1 OAI21X1_5454 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(_14545__bF_buf2), .C(_14619_), .Y(_14620_) );
	INVX1 INVX1_2117 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_17_), .Y(_14621_) );
	OAI21X1 OAI21X1_5455 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14621_), .C(_14558_), .Y(_14622_) );
	OAI21X1 OAI21X1_5456 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(biu_ins_28_bF_buf3), .C(_14622_), .Y(_14623_) );
	XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_14620_), .B(_14623_), .Y(_14624_) );
	XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_14624_), .Y(_14625_) );
	OAI21X1 OAI21X1_5457 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_17_), .B(_14324__bF_buf1), .C(_14328__bF_buf0), .Y(_14626_) );
	AOI21X1 AOI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_14625_), .B(_14324__bF_buf0), .C(_14626_), .Y(_13986__17_) );
	INVX1 INVX1_2118 ( .gnd(gnd), .vdd(vdd), .A(_14620_), .Y(_14627_) );
	NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_14623_), .B(_14627_), .Y(_14628_) );
	OAI21X1 OAI21X1_5458 ( .gnd(gnd), .vdd(vdd), .A(_14627_), .B(_14623_), .C(_14614_), .Y(_14629_) );
	NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_14628_), .B(_14629_), .Y(_14630_) );
	AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_14471_), .B(_14599_), .Y(_14631_) );
	NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_14624_), .B(_14615_), .Y(_14632_) );
	OAI21X1 OAI21X1_5459 ( .gnd(gnd), .vdd(vdd), .A(_14605_), .B(_14631_), .C(_14632_), .Y(_14633_) );
	AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_14633_), .B(_14630_), .Y(_14634_) );
	AOI22X1 AOI22X1_702 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(biu_pc_18_), .C(csr_gpr_iu_rs1_18_), .D(_14334__bF_buf2), .Y(_14635_) );
	OAI21X1 OAI21X1_5460 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(_14545__bF_buf1), .C(_14635_), .Y(_14636_) );
	INVX1 INVX1_2119 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_18_), .Y(_14637_) );
	OAI21X1 OAI21X1_5461 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14637_), .C(_14558_), .Y(_14638_) );
	OAI21X1 OAI21X1_5462 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(biu_ins_29_bF_buf1), .C(_14638_), .Y(_14639_) );
	XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_14636_), .B(_14639_), .Y(_14640_) );
	INVX1 INVX1_2120 ( .gnd(gnd), .vdd(vdd), .A(_14640_), .Y(_14641_) );
	XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_14634_), .B(_14641_), .Y(_14642_) );
	OAI21X1 OAI21X1_5463 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_18_), .B(_14324__bF_buf8), .C(_14328__bF_buf5), .Y(_14643_) );
	AOI21X1 AOI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_14642_), .B(_14324__bF_buf7), .C(_14643_), .Y(_13986__18_) );
	INVX1 INVX1_2121 ( .gnd(gnd), .vdd(vdd), .A(_14636_), .Y(_14644_) );
	NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_14639_), .B(_14644_), .Y(_14645_) );
	INVX1 INVX1_2122 ( .gnd(gnd), .vdd(vdd), .A(_14645_), .Y(_14646_) );
	OAI21X1 OAI21X1_5464 ( .gnd(gnd), .vdd(vdd), .A(_14641_), .B(_14634_), .C(_14646_), .Y(_14647_) );
	AOI22X1 AOI22X1_703 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(biu_pc_19_), .C(csr_gpr_iu_rs1_19_), .D(_14334__bF_buf1), .Y(_14648_) );
	OAI21X1 OAI21X1_5465 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(_14545__bF_buf0), .C(_14648_), .Y(_14649_) );
	INVX1 INVX1_2123 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_19_), .Y(_14650_) );
	OAI21X1 OAI21X1_5466 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(_14650_), .C(_14558_), .Y(_14651_) );
	OAI21X1 OAI21X1_5467 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(biu_ins_30_bF_buf2), .C(_14651_), .Y(_14652_) );
	INVX1 INVX1_2124 ( .gnd(gnd), .vdd(vdd), .A(_14652_), .Y(_14653_) );
	NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .B(_14653_), .Y(_14654_) );
	OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_14653_), .B(_14649_), .Y(_14655_) );
	NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_14654_), .B(_14655_), .Y(_14656_) );
	XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_14647_), .B(_14656_), .Y(_14657_) );
	OAI21X1 OAI21X1_5468 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_19_), .B(_14324__bF_buf6), .C(_14328__bF_buf4), .Y(_14658_) );
	AOI21X1 AOI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_14657_), .B(_14324__bF_buf5), .C(_14658_), .Y(_13986__19_) );
	NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14654_), .B(_14655_), .C(_14640_), .Y(_14659_) );
	OAI21X1 OAI21X1_5469 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .B(_14653_), .C(_14645_), .Y(_14660_) );
	AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_14660_), .B(_14654_), .Y(_14661_) );
	OAI21X1 OAI21X1_5470 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .B(_14630_), .C(_14661_), .Y(_14662_) );
	INVX1 INVX1_2125 ( .gnd(gnd), .vdd(vdd), .A(_14662_), .Y(_14663_) );
	INVX1 INVX1_2126 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .Y(_14664_) );
	NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_14632_), .B(_14664_), .Y(_14665_) );
	OAI21X1 OAI21X1_5471 ( .gnd(gnd), .vdd(vdd), .A(_14665_), .B(_14606_), .C(_14663_), .Y(_14666_) );
	INVX1 INVX1_2127 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_20_), .Y(_14667_) );
	AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(biu_ins_31_bF_buf0), .Y(_14668_) );
	AOI21X1 AOI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_14557_), .B(_14325_), .C(_14668_), .Y(_14669_) );
	OAI21X1 OAI21X1_5472 ( .gnd(gnd), .vdd(vdd), .A(_14667_), .B(_14332_), .C(_14669_), .Y(_14670_) );
	AOI22X1 AOI22X1_704 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_pc_20_), .C(csr_gpr_iu_rs1_20_), .D(_14334__bF_buf0), .Y(_14671_) );
	OAI21X1 OAI21X1_5473 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(_14545__bF_buf3), .C(_14671_), .Y(_14672_) );
	XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14672_), .B(_14670_), .Y(_14673_) );
	XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_14666_), .B(_14673_), .Y(_14674_) );
	OAI21X1 OAI21X1_5474 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_20_), .B(_14324__bF_buf4), .C(_14328__bF_buf3), .Y(_14675_) );
	AOI21X1 AOI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_14674_), .B(_14324__bF_buf3), .C(_14675_), .Y(_13986__20_) );
	NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_14670_), .B(_14672_), .Y(_14676_) );
	NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_14673_), .B(_14666_), .Y(_14677_) );
	NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_14676_), .B(_14677_), .Y(_14678_) );
	INVX1 INVX1_2128 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_21_), .Y(_14679_) );
	OAI21X1 OAI21X1_5475 ( .gnd(gnd), .vdd(vdd), .A(_14679_), .B(_14332_), .C(_14669_), .Y(_14680_) );
	AOI22X1 AOI22X1_705 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_pc_21_), .C(csr_gpr_iu_rs1_21_), .D(_14334__bF_buf4), .Y(_14681_) );
	OAI21X1 OAI21X1_5476 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(_14545__bF_buf2), .C(_14681_), .Y(_14682_) );
	XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_14682_), .B(_14680_), .Y(_14683_) );
	XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_14678_), .B(_14683_), .Y(_14684_) );
	OAI21X1 OAI21X1_5477 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_21_), .B(_14324__bF_buf2), .C(_14328__bF_buf2), .Y(_14685_) );
	AOI21X1 AOI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .B(_14324__bF_buf1), .C(_14685_), .Y(_13986__21_) );
	NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_14680_), .B(_14682_), .Y(_14686_) );
	NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_14676_), .B(_14686_), .Y(_14687_) );
	NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_14673_), .B(_14683_), .Y(_14688_) );
	INVX1 INVX1_2129 ( .gnd(gnd), .vdd(vdd), .A(_14688_), .Y(_14689_) );
	AOI21X1 AOI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_14666_), .B(_14689_), .C(_14687_), .Y(_14690_) );
	INVX1 INVX1_2130 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_22_), .Y(_14691_) );
	OAI21X1 OAI21X1_5478 ( .gnd(gnd), .vdd(vdd), .A(_14691_), .B(_14332_), .C(_14669_), .Y(_14692_) );
	AOI22X1 AOI22X1_706 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_pc_22_), .C(csr_gpr_iu_rs1_22_), .D(_14334__bF_buf3), .Y(_14693_) );
	OAI21X1 OAI21X1_5479 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(_14545__bF_buf1), .C(_14693_), .Y(_14694_) );
	NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_14692_), .B(_14694_), .Y(_14695_) );
	NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_14692_), .B(_14694_), .Y(_14696_) );
	INVX1 INVX1_2131 ( .gnd(gnd), .vdd(vdd), .A(_14696_), .Y(_14697_) );
	NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_14695_), .B(_14697_), .Y(_14698_) );
	INVX1 INVX1_2132 ( .gnd(gnd), .vdd(vdd), .A(_14698_), .Y(_14699_) );
	XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_14690_), .B(_14699_), .Y(_14700_) );
	OAI21X1 OAI21X1_5480 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_22_), .B(_14324__bF_buf0), .C(_14328__bF_buf1), .Y(_14701_) );
	AOI21X1 AOI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_14700_), .B(_14324__bF_buf8), .C(_14701_), .Y(_13986__22_) );
	OAI21X1 OAI21X1_5481 ( .gnd(gnd), .vdd(vdd), .A(_14699_), .B(_14690_), .C(_14696_), .Y(_14702_) );
	INVX1 INVX1_2133 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_23_), .Y(_14703_) );
	OAI21X1 OAI21X1_5482 ( .gnd(gnd), .vdd(vdd), .A(_14703_), .B(_14332_), .C(_14669_), .Y(_14704_) );
	AOI22X1 AOI22X1_707 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(biu_pc_23_), .C(csr_gpr_iu_rs1_23_), .D(_14334__bF_buf2), .Y(_14705_) );
	OAI21X1 OAI21X1_5483 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(_14545__bF_buf0), .C(_14705_), .Y(_14706_) );
	NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14706_), .Y(_14707_) );
	NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14706_), .Y(_14708_) );
	INVX1 INVX1_2134 ( .gnd(gnd), .vdd(vdd), .A(_14708_), .Y(_14709_) );
	NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_14707_), .B(_14709_), .Y(_14710_) );
	XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_14702_), .B(_14710_), .Y(_14711_) );
	OAI21X1 OAI21X1_5484 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_23_), .B(_14324__bF_buf7), .C(_14328__bF_buf0), .Y(_14712_) );
	AOI21X1 AOI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_14711_), .B(_14324__bF_buf6), .C(_14712_), .Y(_13986__23_) );
	NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_14698_), .B(_14710_), .Y(_14713_) );
	NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_14688_), .B(_14713_), .Y(_14714_) );
	NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(_14632_), .B(_14664_), .C(_14714_), .Y(_14715_) );
	NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(_14687_), .B(_14698_), .C(_14710_), .Y(_14716_) );
	NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(_14696_), .B(_14708_), .C(_14716_), .Y(_14717_) );
	AOI21X1 AOI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_14662_), .B(_14714_), .C(_14717_), .Y(_14718_) );
	OAI21X1 OAI21X1_5485 ( .gnd(gnd), .vdd(vdd), .A(_14715_), .B(_14606_), .C(_14718_), .Y(_14719_) );
	INVX1 INVX1_2135 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_24_), .Y(_14720_) );
	OAI21X1 OAI21X1_5486 ( .gnd(gnd), .vdd(vdd), .A(_14720_), .B(_14332_), .C(_14669_), .Y(_14721_) );
	AOI22X1 AOI22X1_708 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_pc_24_), .C(csr_gpr_iu_rs1_24_), .D(_14334__bF_buf1), .Y(_14722_) );
	OAI21X1 OAI21X1_5487 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(_14545__bF_buf3), .C(_14722_), .Y(_14723_) );
	NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_14721_), .B(_14723_), .Y(_14724_) );
	INVX2 INVX2_193 ( .gnd(gnd), .vdd(vdd), .A(_14724_), .Y(_14725_) );
	NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_14721_), .B(_14723_), .Y(_14726_) );
	NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_14726_), .B(_14725_), .Y(_14727_) );
	NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_14727_), .B(_14719_), .Y(_14728_) );
	INVX1 INVX1_2136 ( .gnd(gnd), .vdd(vdd), .A(_14719_), .Y(_14729_) );
	OAI21X1 OAI21X1_5488 ( .gnd(gnd), .vdd(vdd), .A(_14725_), .B(_14726_), .C(_14729_), .Y(_14730_) );
	NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_14728_), .B(_14730_), .Y(_14731_) );
	OAI21X1 OAI21X1_5489 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_24_), .B(_14324__bF_buf5), .C(_14328__bF_buf5), .Y(_14732_) );
	AOI21X1 AOI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_14731_), .B(_14324__bF_buf4), .C(_14732_), .Y(_13986__24_) );
	OAI21X1 OAI21X1_5490 ( .gnd(gnd), .vdd(vdd), .A(_14726_), .B(_14729_), .C(_14724_), .Y(_14733_) );
	INVX1 INVX1_2137 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_25_), .Y(_14734_) );
	OAI21X1 OAI21X1_5491 ( .gnd(gnd), .vdd(vdd), .A(_14734_), .B(_14332_), .C(_14669_), .Y(_14735_) );
	AOI22X1 AOI22X1_709 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_pc_25_), .C(csr_gpr_iu_rs1_25_), .D(_14334__bF_buf0), .Y(_14736_) );
	OAI21X1 OAI21X1_5492 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(_14545__bF_buf2), .C(_14736_), .Y(_14737_) );
	NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_14735_), .B(_14737_), .Y(_14738_) );
	INVX1 INVX1_2138 ( .gnd(gnd), .vdd(vdd), .A(_14738_), .Y(_14739_) );
	NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_14735_), .B(_14737_), .Y(_14740_) );
	NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_14740_), .B(_14739_), .Y(_14741_) );
	XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_14733_), .B(_14741_), .Y(_14742_) );
	OAI21X1 OAI21X1_5493 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_25_), .B(_14324__bF_buf3), .C(_14328__bF_buf4), .Y(_14743_) );
	AOI21X1 AOI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_14742_), .B(_14324__bF_buf2), .C(_14743_), .Y(_13986__25_) );
	NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_14727_), .B(_14741_), .Y(_14744_) );
	INVX1 INVX1_2139 ( .gnd(gnd), .vdd(vdd), .A(_14744_), .Y(_14745_) );
	NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_14725_), .B(_14739_), .Y(_14746_) );
	INVX1 INVX1_2140 ( .gnd(gnd), .vdd(vdd), .A(_14746_), .Y(_14747_) );
	AOI21X1 AOI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_14719_), .B(_14745_), .C(_14747_), .Y(_14748_) );
	INVX1 INVX1_2141 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_26_), .Y(_14749_) );
	OAI21X1 OAI21X1_5494 ( .gnd(gnd), .vdd(vdd), .A(_14749_), .B(_14332_), .C(_14669_), .Y(_14750_) );
	AOI22X1 AOI22X1_710 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_pc_26_), .C(csr_gpr_iu_rs1_26_), .D(_14334__bF_buf4), .Y(_14751_) );
	OAI21X1 OAI21X1_5495 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(_14545__bF_buf1), .C(_14751_), .Y(_14752_) );
	XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_14752_), .B(_14750_), .Y(_14753_) );
	XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_14748_), .B(_14753_), .Y(_14754_) );
	OAI21X1 OAI21X1_5496 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_26_), .B(_14324__bF_buf1), .C(_14328__bF_buf3), .Y(_14755_) );
	AOI21X1 AOI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_14754_), .B(_14324__bF_buf0), .C(_14755_), .Y(_13986__26_) );
	NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_14750_), .B(_14752_), .Y(_14756_) );
	OAI21X1 OAI21X1_5497 ( .gnd(gnd), .vdd(vdd), .A(_14753_), .B(_14748_), .C(_14756_), .Y(_14757_) );
	INVX1 INVX1_2142 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_27_), .Y(_14758_) );
	OAI21X1 OAI21X1_5498 ( .gnd(gnd), .vdd(vdd), .A(_14758_), .B(_14332_), .C(_14669_), .Y(_14759_) );
	AOI22X1 AOI22X1_711 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf4), .B(biu_pc_27_), .C(csr_gpr_iu_rs1_27_), .D(_14334__bF_buf3), .Y(_14760_) );
	OAI21X1 OAI21X1_5499 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(_14545__bF_buf0), .C(_14760_), .Y(_14761_) );
	XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_14761_), .B(_14759_), .Y(_14762_) );
	XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14757_), .B(_14762_), .Y(_14763_) );
	OAI21X1 OAI21X1_5500 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_27_), .B(_14324__bF_buf8), .C(_14328__bF_buf2), .Y(_14764_) );
	AOI21X1 AOI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_14763_), .B(_14324__bF_buf7), .C(_14764_), .Y(_13986__27_) );
	NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_14753_), .B(_14762_), .Y(_14765_) );
	AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_14745_), .B(_14765_), .Y(_14766_) );
	OAI21X1 OAI21X1_5501 ( .gnd(gnd), .vdd(vdd), .A(_14725_), .B(_14739_), .C(_14765_), .Y(_14767_) );
	AOI22X1 AOI22X1_712 ( .gnd(gnd), .vdd(vdd), .A(_14752_), .B(_14750_), .C(_14759_), .D(_14761_), .Y(_14768_) );
	NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_14768_), .B(_14767_), .Y(_14769_) );
	AOI21X1 AOI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_14719_), .B(_14766_), .C(_14769_), .Y(_14770_) );
	INVX1 INVX1_2143 ( .gnd(gnd), .vdd(vdd), .A(_14669_), .Y(_14771_) );
	AOI21X1 AOI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_28_), .B(_14331__bF_buf3), .C(_14771_), .Y(_14772_) );
	INVX1 INVX1_2144 ( .gnd(gnd), .vdd(vdd), .A(_14772_), .Y(_14773_) );
	AOI22X1 AOI22X1_713 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf2), .B(biu_pc_28_), .C(csr_gpr_iu_rs1_28_), .D(_14334__bF_buf2), .Y(_14774_) );
	OAI21X1 OAI21X1_5502 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf1), .B(_14545__bF_buf3), .C(_14774_), .Y(_14775_) );
	NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_14775_), .B(_14773_), .Y(_14776_) );
	NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_14775_), .B(_14773_), .Y(_14777_) );
	INVX1 INVX1_2145 ( .gnd(gnd), .vdd(vdd), .A(_14777_), .Y(_14778_) );
	NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_14776_), .B(_14778_), .Y(_14779_) );
	XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .B(_14779_), .Y(_14780_) );
	OAI21X1 OAI21X1_5503 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_28_), .B(_14324__bF_buf6), .C(_14328__bF_buf1), .Y(_14781_) );
	AOI21X1 AOI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_14780_), .B(_14324__bF_buf5), .C(_14781_), .Y(_13986__28_) );
	INVX1 INVX1_2146 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .Y(_14782_) );
	AOI21X1 AOI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_14782_), .B(_14779_), .C(_14778_), .Y(_14783_) );
	AOI21X1 AOI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_29_), .B(_14331__bF_buf2), .C(_14771_), .Y(_14784_) );
	AOI22X1 AOI22X1_714 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf0), .B(biu_pc_29_), .C(csr_gpr_iu_rs1_29_), .D(_14334__bF_buf1), .Y(_14785_) );
	OAI21X1 OAI21X1_5504 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf7), .B(_14545__bF_buf2), .C(_14785_), .Y(_14786_) );
	XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_14784_), .B(_14786_), .Y(_14787_) );
	OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_14783_), .B(_14787_), .Y(_14788_) );
	INVX8 INVX8_106 ( .gnd(gnd), .vdd(vdd), .A(_14324__bF_buf4), .Y(_14789_) );
	AOI21X1 AOI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_14783_), .B(_14787_), .C(_14789__bF_buf4), .Y(_14790_) );
	OAI21X1 OAI21X1_5505 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_29_), .B(_14324__bF_buf3), .C(_14328__bF_buf0), .Y(_14791_) );
	AOI21X1 AOI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_14788_), .B(_14790_), .C(_14791_), .Y(_13986__29_) );
	NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_14787_), .B(_14779_), .Y(_14792_) );
	INVX1 INVX1_2147 ( .gnd(gnd), .vdd(vdd), .A(_14784_), .Y(_14793_) );
	AOI21X1 AOI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_14793_), .B(_14786_), .C(_14778_), .Y(_14794_) );
	OAI21X1 OAI21X1_5506 ( .gnd(gnd), .vdd(vdd), .A(_14792_), .B(_14770_), .C(_14794_), .Y(_14795_) );
	AOI21X1 AOI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_30_), .B(_14331__bF_buf1), .C(_14771_), .Y(_14796_) );
	AOI22X1 AOI22X1_715 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf6), .B(biu_pc_30_), .C(csr_gpr_iu_rs1_30_), .D(_14334__bF_buf0), .Y(_14797_) );
	OAI21X1 OAI21X1_5507 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf5), .B(_14545__bF_buf1), .C(_14797_), .Y(_14798_) );
	XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_14796_), .B(_14798_), .Y(_14799_) );
	XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_14795_), .B(_14799_), .Y(_14800_) );
	OAI21X1 OAI21X1_5508 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_30_), .B(_14324__bF_buf2), .C(_14328__bF_buf5), .Y(_14801_) );
	AOI21X1 AOI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_14800_), .B(_14324__bF_buf1), .C(_14801_), .Y(_13986__30_) );
	AOI21X1 AOI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_14535_), .B(_14797_), .C(_14796_), .Y(_14802_) );
	AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_14795_), .B(_14799_), .Y(_14803_) );
	INVX1 INVX1_2148 ( .gnd(gnd), .vdd(vdd), .A(biu_pc_31_), .Y(_14804_) );
	OAI21X1 OAI21X1_5509 ( .gnd(gnd), .vdd(vdd), .A(_14804_), .B(_14332_), .C(_14669_), .Y(_14805_) );
	AOI21X1 AOI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jalr), .B(csr_gpr_iu_rs1_31_), .C(csr_gpr_iu_ins_dec_jal_bF_buf4), .Y(_14806_) );
	AOI22X1 AOI22X1_716 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_jal_bF_buf3), .B(_14804_), .C(_14806_), .D(_14545__bF_buf0), .Y(_14807_) );
	XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14807_), .B(_14805_), .Y(_14808_) );
	INVX1 INVX1_2149 ( .gnd(gnd), .vdd(vdd), .A(_14808_), .Y(_14809_) );
	OAI21X1 OAI21X1_5510 ( .gnd(gnd), .vdd(vdd), .A(_14802_), .B(_14803_), .C(_14809_), .Y(_14810_) );
	AOI21X1 AOI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_14795_), .B(_14799_), .C(_14802_), .Y(_14811_) );
	AOI21X1 AOI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_14811_), .B(_14808_), .C(_14789__bF_buf3), .Y(_14812_) );
	OAI21X1 OAI21X1_5511 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csr_pc_next_31_), .B(_14324__bF_buf0), .C(_14328__bF_buf4), .Y(_14813_) );
	AOI21X1 AOI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_14812_), .B(_14810_), .C(_14813_), .Y(_13986__31_) );
	NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(amoxor_bF_buf1), .B(csr_gpr_iu_ins_dec_sc_w), .Y(_14814_) );
	NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(amomax), .B(amomaxu), .Y(_14815_) );
	NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_14814_), .B(_14815_), .Y(_14816_) );
	OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_ins_dec_lr_w), .B(amoadd_bF_buf0), .Y(_14817_) );
	NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(amoswap), .B(_14817_), .Y(_14818_) );
	NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(amomin), .B(amoor), .Y(_14819_) );
	NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(amominu), .B(amoand), .Y(_14820_) );
	NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(_14819_), .B(_14820_), .C(_14818_), .Y(_14821_) );
	NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_14816_), .B(_14821_), .Y(_14822_) );
	INVX1 INVX1_2150 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .Y(_14823_) );
	NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(biu_exce_chk_opc_0_), .Y(_14824_) );
	INVX8 INVX8_107 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .Y(_14825_) );
	AOI21X1 AOI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_14823_), .B(csr_gpr_iu_csrrw), .C(_14825__bF_buf4), .Y(_14826_) );
	INVX1 INVX1_2151 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_18_), .Y(_14827_) );
	INVX1 INVX1_2152 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_19_), .Y(_14828_) );
	NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_16_), .B(csr_gpr_iu_rs1_17_), .Y(_14829_) );
	NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(_14827_), .B(_14828_), .C(_14829_), .Y(_14830_) );
	INVX1 INVX1_2153 ( .gnd(gnd), .vdd(vdd), .A(_14830_), .Y(_14831_) );
	NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_20_), .B(csr_gpr_iu_rs1_21_), .Y(_14832_) );
	NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_22_), .B(csr_gpr_iu_rs1_23_), .Y(_14833_) );
	NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_14832_), .B(_14833_), .Y(_14834_) );
	INVX1 INVX1_2154 ( .gnd(gnd), .vdd(vdd), .A(_14834_), .Y(_14835_) );
	INVX1 INVX1_2155 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_14_), .Y(_14836_) );
	INVX1 INVX1_2156 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_15_), .Y(_14837_) );
	NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .B(csr_gpr_iu_rs1_13_), .Y(_14838_) );
	NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(_14836_), .B(_14837_), .C(_14838_), .Y(_14839_) );
	INVX1 INVX1_2157 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_24_), .Y(_14840_) );
	INVX1 INVX1_2158 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_25_), .Y(_14841_) );
	NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_26_), .B(csr_gpr_iu_rs1_27_), .Y(_14842_) );
	NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(_14840_), .B(_14841_), .C(_14842_), .Y(_14843_) );
	NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_14839_), .B(_14843_), .Y(_14844_) );
	NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(_14831_), .B(_14835_), .C(_14844_), .Y(_14845_) );
	INVX1 INVX1_2159 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .Y(_14846_) );
	INVX1 INVX1_2160 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_11_), .Y(_14847_) );
	NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_30_), .B(csr_gpr_iu_rs1_31_), .Y(_14848_) );
	NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(_14846_), .B(_14847_), .C(_14848_), .Y(_14849_) );
	INVX1 INVX1_2161 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .Y(_14850_) );
	INVX1 INVX1_2162 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_7_), .Y(_14851_) );
	NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .B(csr_gpr_iu_rs1_9_), .Y(_14852_) );
	NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(_14850_), .B(_14851_), .C(_14852_), .Y(_14853_) );
	NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_14849_), .B(_14853_), .Y(_14854_) );
	INVX1 INVX1_2163 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_4_), .Y(_14855_) );
	INVX1 INVX1_2164 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .Y(_14856_) );
	NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .B(csr_gpr_iu_rs1_3_), .Y(_14857_) );
	NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(_14855_), .B(_14856_), .C(_14857_), .Y(_14858_) );
	INVX1 INVX1_2165 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_1_), .Y(_14859_) );
	NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_28_), .B(csr_gpr_iu_rs1_29_), .Y(_14860_) );
	NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(_14823_), .B(_14859_), .C(_14860_), .Y(_14861_) );
	NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_14858_), .B(_14861_), .Y(_14862_) );
	NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_14854_), .B(_14862_), .Y(_14863_) );
	INVX1 INVX1_2166 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrc), .Y(_14864_) );
	NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(csr_0_), .B(_14864_), .Y(_14865_) );
	OAI21X1 OAI21X1_5512 ( .gnd(gnd), .vdd(vdd), .A(_14863_), .B(_14845_), .C(_14865_), .Y(_14866_) );
	INVX1 INVX1_2167 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_15_bF_buf2), .Y(_14867_) );
	NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrsi), .B(csr_gpr_iu_csrrwi), .Y(_14868_) );
	INVX1 INVX1_2168 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrwi), .Y(_14869_) );
	AOI21X1 AOI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(csr_0_), .B(_14869_), .C(_14868_), .Y(_14870_) );
	OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_16_), .B(biu_ins_15_bF_buf1), .Y(_14871_) );
	INVX1 INVX1_2169 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_19_), .Y(_14872_) );
	NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .B(biu_ins_17_), .Y(_14873_) );
	NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_14872_), .B(_14873_), .Y(_14874_) );
	NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_14871_), .B(_14874_), .Y(_14875_) );
	OAI21X1 OAI21X1_5513 ( .gnd(gnd), .vdd(vdd), .A(csr_0_), .B(_14875_), .C(csr_gpr_iu_csrrci), .Y(_14876_) );
	AOI22X1 AOI22X1_717 ( .gnd(gnd), .vdd(vdd), .A(_14867_), .B(_14870_), .C(_14868_), .D(_14876_), .Y(_14877_) );
	OAI21X1 OAI21X1_5514 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrc), .B(_14877_), .C(_14866_), .Y(_14878_) );
	OAI21X1 OAI21X1_5515 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .B(csr_0_), .C(csr_gpr_iu_csrrs), .Y(_14879_) );
	OAI21X1 OAI21X1_5516 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrs), .B(_14878_), .C(_14879_), .Y(_14880_) );
	OAI21X1 OAI21X1_5517 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrw), .B(_14880_), .C(_14826_), .Y(_14881_) );
	AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .B(csr_gpr_iu_imm12_0_), .Y(_14882_) );
	NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf4), .B(_14882_), .Y(_14883_) );
	OAI21X1 OAI21X1_5518 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .B(csr_gpr_iu_imm12_0_), .C(_14883_), .Y(_14884_) );
	NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(_14822__bF_buf3), .B(_14884_), .C(_14881_), .Y(_14885_) );
	OAI21X1 OAI21X1_5519 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_0_), .B(_14822__bF_buf2), .C(_14885_), .Y(_14886_) );
	OAI21X1 OAI21X1_5520 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_0_), .B(_14324__bF_buf8), .C(_14328__bF_buf3), .Y(_14887_) );
	AOI21X1 AOI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .B(_14324__bF_buf7), .C(_14887_), .Y(_13985__0_) );
	XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_1_), .B(csr_gpr_iu_imm12_1_), .Y(_14888_) );
	NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .B(_14888_), .Y(_14889_) );
	NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .B(_14888_), .Y(_14890_) );
	OAI21X1 OAI21X1_5521 ( .gnd(gnd), .vdd(vdd), .A(biu_exce_chk_opc_1_), .B(biu_exce_chk_opc_0_), .C(_14890_), .Y(_14891_) );
	NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14891_), .Y(_14892_) );
	NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrs), .B(csr_gpr_iu_csrrw), .Y(_14893_) );
	NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrci), .B(csr_gpr_iu_csrrsi), .Y(_14894_) );
	NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrc), .B(csr_gpr_iu_csrrs), .Y(_14895_) );
	OAI21X1 OAI21X1_5522 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrwi), .B(_14894_), .C(_14895_), .Y(_14896_) );
	OAI21X1 OAI21X1_5523 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrsi), .B(csr_gpr_iu_csrrwi), .C(_14895_), .Y(_14897_) );
	INVX1 INVX1_2170 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14898_) );
	AOI22X1 AOI22X1_718 ( .gnd(gnd), .vdd(vdd), .A(csr_1_), .B(_14896__bF_buf4), .C(biu_ins_16_), .D(_14898_), .Y(_14899_) );
	OAI22X1 OAI22X1_834 ( .gnd(gnd), .vdd(vdd), .A(_14859_), .B(_14893_), .C(csr_gpr_iu_csrrw), .D(_14899_), .Y(_14900_) );
	AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_14900_), .B(_14824__bF_buf3), .Y(_14901_) );
	OAI21X1 OAI21X1_5524 ( .gnd(gnd), .vdd(vdd), .A(_14892_), .B(_14901_), .C(_14822__bF_buf1), .Y(_14902_) );
	INVX8 INVX8_108 ( .gnd(gnd), .vdd(vdd), .A(_14822__bF_buf0), .Y(_14903_) );
	AOI21X1 AOI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(csr_gpr_iu_rs1_1_), .C(_14789__bF_buf2), .Y(_14904_) );
	OAI21X1 OAI21X1_5525 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_1_), .B(_14324__bF_buf6), .C(_14328__bF_buf2), .Y(_14905_) );
	AOI21X1 AOI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .B(_14904_), .C(_14905_), .Y(_13985__1_) );
	OAI21X1 OAI21X1_5526 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf2), .B(_14323__bF_buf2), .C(addr_csr_2_), .Y(_14906_) );
	OAI21X1 OAI21X1_5527 ( .gnd(gnd), .vdd(vdd), .A(_14859_), .B(_14349_), .C(_14890_), .Y(_14907_) );
	NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(_14371_), .Y(_14908_) );
	NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_2_), .B(csr_gpr_iu_imm12_2_), .Y(_14909_) );
	NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_14909_), .B(_14908_), .Y(_14910_) );
	XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_14907_), .B(_14910_), .Y(_14911_) );
	INVX8 INVX8_109 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrw), .Y(_14912_) );
	AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_14896__bF_buf3), .B(csr_2_), .Y(_14913_) );
	AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .B(biu_ins_17_), .Y(_14914_) );
	OAI21X1 OAI21X1_5528 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .B(_14914_), .C(_14912__bF_buf4), .Y(_14915_) );
	INVX8 INVX8_110 ( .gnd(gnd), .vdd(vdd), .A(_14893_), .Y(_14916_) );
	AOI21X1 AOI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_14916__bF_buf3), .B(csr_gpr_iu_rs1_2_), .C(_14825__bF_buf3), .Y(_14917_) );
	AOI22X1 AOI22X1_719 ( .gnd(gnd), .vdd(vdd), .A(_14915_), .B(_14917_), .C(_14825__bF_buf2), .D(_14911_), .Y(_14918_) );
	AOI21X1 AOI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_14357_), .C(_14789__bF_buf1), .Y(_14919_) );
	OAI21X1 OAI21X1_5529 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14918_), .C(_14919_), .Y(_14920_) );
	AOI21X1 AOI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .B(_14906_), .C(rst_bF_buf48), .Y(_13985__2_) );
	OAI21X1 OAI21X1_5530 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf1), .B(_14323__bF_buf1), .C(addr_csr_3_), .Y(_14921_) );
	NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_14910_), .B(_14907_), .Y(_14922_) );
	OAI21X1 OAI21X1_5531 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(_14371_), .C(_14922_), .Y(_14923_) );
	NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .B(csr_gpr_iu_imm12_3_), .Y(_14924_) );
	INVX1 INVX1_2171 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_3_), .Y(_14925_) );
	NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_14925_), .B(_14385_), .Y(_14926_) );
	NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .B(_14926_), .Y(_14927_) );
	AOI21X1 AOI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_14923_), .B(_14927_), .C(_14824__bF_buf2), .Y(_14928_) );
	OAI21X1 OAI21X1_5532 ( .gnd(gnd), .vdd(vdd), .A(_14923_), .B(_14927_), .C(_14928_), .Y(_14929_) );
	INVX1 INVX1_2172 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_18_), .Y(_14930_) );
	NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(csr_3_), .B(_14896__bF_buf2), .Y(_14931_) );
	OAI21X1 OAI21X1_5533 ( .gnd(gnd), .vdd(vdd), .A(_14930_), .B(_14897_), .C(_14931_), .Y(_14932_) );
	NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(_14824__bF_buf1), .C(_14932_), .Y(_14933_) );
	AOI21X1 AOI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_14929_), .B(_14933_), .C(_14903__bF_buf2), .Y(_14934_) );
	OAI21X1 OAI21X1_5534 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrs), .B(csr_gpr_iu_csrrw), .C(_14824__bF_buf0), .Y(_14935_) );
	AOI21X1 AOI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_14822__bF_buf3), .B(_14935_), .C(_14925_), .Y(_14936_) );
	OAI21X1 OAI21X1_5535 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .B(_14934_), .C(_14324__bF_buf5), .Y(_14937_) );
	AOI21X1 AOI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_14937_), .B(_14921_), .C(rst_bF_buf47), .Y(_13985__3_) );
	OAI21X1 OAI21X1_5536 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf0), .B(_14323__bF_buf0), .C(addr_csr_4_), .Y(_14938_) );
	AOI21X1 AOI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_14822__bF_buf2), .B(_14935_), .C(_14855_), .Y(_14939_) );
	NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_4_), .B(csr_gpr_iu_imm12_4_), .Y(_14940_) );
	NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_14855_), .B(_14404_), .Y(_14941_) );
	NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14941_), .Y(_14942_) );
	AOI21X1 AOI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_14927_), .B(_14908_), .C(_14926_), .Y(_14943_) );
	NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(_14910_), .B(_14927_), .C(_14907_), .Y(_14944_) );
	NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_14943_), .B(_14944_), .Y(_14945_) );
	AOI21X1 AOI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_14942_), .C(_14824__bF_buf5), .Y(_14946_) );
	OAI21X1 OAI21X1_5537 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .B(_14945_), .C(_14946_), .Y(_14947_) );
	NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(csr_4_), .B(_14896__bF_buf1), .Y(_14948_) );
	OAI21X1 OAI21X1_5538 ( .gnd(gnd), .vdd(vdd), .A(_14872_), .B(_14897_), .C(_14948_), .Y(_14949_) );
	NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf2), .B(_14824__bF_buf4), .C(_14949_), .Y(_14950_) );
	AOI21X1 AOI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14950_), .C(_14903__bF_buf1), .Y(_14951_) );
	OAI21X1 OAI21X1_5539 ( .gnd(gnd), .vdd(vdd), .A(_14939_), .B(_14951_), .C(_14324__bF_buf4), .Y(_14952_) );
	AOI21X1 AOI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .B(_14938_), .C(rst_bF_buf46), .Y(_13985__4_) );
	OAI21X1 OAI21X1_5540 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf3), .B(_14323__bF_buf3), .C(addr_csr_5_), .Y(_14953_) );
	INVX1 INVX1_2173 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .Y(_14954_) );
	INVX1 INVX1_2174 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .Y(_14955_) );
	OAI21X1 OAI21X1_5541 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14955_), .C(_14954_), .Y(_14956_) );
	NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .B(biu_ins_25_bF_buf0), .Y(_14957_) );
	NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_14856_), .B(_14425_), .Y(_14958_) );
	NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_14957_), .B(_14958_), .Y(_14959_) );
	OAI21X1 OAI21X1_5542 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14956_), .C(_14825__bF_buf1), .Y(_14960_) );
	AOI21X1 AOI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_14959_), .C(_14960_), .Y(_14961_) );
	AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf1), .B(csr_5_), .Y(_14962_) );
	AOI22X1 AOI22X1_720 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_5_), .B(_14916__bF_buf2), .C(_14962_), .D(_14896__bF_buf0), .Y(_14963_) );
	OAI21X1 OAI21X1_5543 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf0), .B(_14963_), .C(_14822__bF_buf1), .Y(_14964_) );
	AOI21X1 AOI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_14856_), .C(_14789__bF_buf0), .Y(_14965_) );
	OAI21X1 OAI21X1_5544 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_14961_), .C(_14965_), .Y(_14966_) );
	AOI21X1 AOI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_14966_), .B(_14953_), .C(rst_bF_buf45), .Y(_13985__5_) );
	NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .B(_14959_), .Y(_14967_) );
	AOI21X1 AOI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14941_), .C(_14958_), .Y(_14968_) );
	OAI21X1 OAI21X1_5545 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_14955_), .C(_14968_), .Y(_14969_) );
	NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .B(biu_ins_26_bF_buf2), .Y(_14970_) );
	NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_14850_), .B(_14441_), .Y(_14971_) );
	NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_14970_), .B(_14971_), .Y(_14972_) );
	XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_14972_), .Y(_14973_) );
	AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf0), .B(csr_6_), .Y(_14974_) );
	AOI22X1 AOI22X1_721 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_6_), .B(_14916__bF_buf1), .C(_14974_), .D(_14896__bF_buf4), .Y(_14975_) );
	AOI21X1 AOI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf3), .B(_14975_), .C(_14903__bF_buf5), .Y(_14976_) );
	OAI21X1 OAI21X1_5546 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf2), .B(_14973_), .C(_14976_), .Y(_14977_) );
	AOI21X1 AOI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_6_), .C(_14789__bF_buf4), .Y(_14978_) );
	OAI21X1 OAI21X1_5547 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_6_), .B(_14324__bF_buf3), .C(_14328__bF_buf1), .Y(_14979_) );
	AOI21X1 AOI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .B(_14978_), .C(_14979_), .Y(_13985__6_) );
	OAI21X1 OAI21X1_5548 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf2), .B(_14323__bF_buf2), .C(addr_csr_7_), .Y(_14980_) );
	AOI21X1 AOI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_14972_), .C(_14971_), .Y(_14981_) );
	NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_7_), .B(biu_ins_27_bF_buf1), .Y(_14982_) );
	NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_14851_), .B(_14457_), .Y(_14983_) );
	NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14983_), .Y(_14984_) );
	INVX1 INVX1_2175 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_13987_) );
	AOI21X1 AOI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_13987_), .C(_14824__bF_buf1), .Y(_13988_) );
	OAI21X1 OAI21X1_5549 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_13987_), .C(_13988_), .Y(_13989_) );
	INVX2 INVX2_194 ( .gnd(gnd), .vdd(vdd), .A(_14896__bF_buf3), .Y(_13990_) );
	NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(csr_7_), .B(_14912__bF_buf4), .Y(_13991_) );
	OAI22X1 OAI22X1_835 ( .gnd(gnd), .vdd(vdd), .A(_14851_), .B(_14893_), .C(_13991_), .D(_13990_), .Y(_13992_) );
	AOI21X1 AOI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf0), .B(_13992_), .C(_14903__bF_buf3), .Y(_13993_) );
	AOI21X1 AOI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_13989_), .B(_13993_), .C(_14789__bF_buf3), .Y(_13994_) );
	OAI21X1 OAI21X1_5550 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_7_), .B(_14822__bF_buf0), .C(_13994_), .Y(_13995_) );
	AOI21X1 AOI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_13995_), .B(_14980_), .C(rst_bF_buf44), .Y(_13985__7_) );
	AOI21X1 AOI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .B(_14971_), .C(_14983_), .Y(_13996_) );
	NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_14972_), .B(_14984_), .Y(_13997_) );
	OAI21X1 OAI21X1_5551 ( .gnd(gnd), .vdd(vdd), .A(_13997_), .B(_14968_), .C(_13996_), .Y(_13998_) );
	NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_13997_), .Y(_13999_) );
	AOI21X1 AOI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_13999_), .C(_13998_), .Y(_14000_) );
	INVX1 INVX1_2176 ( .gnd(gnd), .vdd(vdd), .A(_14000_), .Y(_14001_) );
	NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .B(biu_ins_28_bF_buf2), .Y(_14002_) );
	INVX1 INVX1_2177 ( .gnd(gnd), .vdd(vdd), .A(_14002_), .Y(_14003_) );
	NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .B(biu_ins_28_bF_buf1), .Y(_14004_) );
	NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_14004_), .B(_14003_), .Y(_14005_) );
	AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_14001_), .B(_14005_), .Y(_14006_) );
	NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_14005_), .B(_14001_), .Y(_14007_) );
	OAI21X1 OAI21X1_5552 ( .gnd(gnd), .vdd(vdd), .A(_14007_), .B(_14006_), .C(_14825__bF_buf4), .Y(_14008_) );
	AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(csr_8_), .Y(_14009_) );
	AOI22X1 AOI22X1_722 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_8_), .B(_14916__bF_buf0), .C(_14009_), .D(_14896__bF_buf2), .Y(_14010_) );
	AOI21X1 AOI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .B(_14010_), .C(_14903__bF_buf2), .Y(_14011_) );
	NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_14011_), .B(_14008_), .Y(_14012_) );
	AOI21X1 AOI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_8_), .C(_14789__bF_buf2), .Y(_14013_) );
	OAI21X1 OAI21X1_5553 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_8_), .B(_14324__bF_buf2), .C(_14328__bF_buf0), .Y(_14014_) );
	AOI21X1 AOI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_14012_), .B(_14013_), .C(_14014_), .Y(_13985__8_) );
	OAI21X1 OAI21X1_5554 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf1), .B(_14323__bF_buf1), .C(addr_csr_9_), .Y(_14015_) );
	OAI21X1 OAI21X1_5555 ( .gnd(gnd), .vdd(vdd), .A(_14004_), .B(_14000_), .C(_14002_), .Y(_14016_) );
	INVX1 INVX1_2178 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_9_), .Y(_14017_) );
	NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_14017_), .B(_14500_), .Y(_14018_) );
	NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_9_), .B(biu_ins_29_bF_buf0), .Y(_14019_) );
	NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_14019_), .B(_14018_), .Y(_14020_) );
	INVX1 INVX1_2179 ( .gnd(gnd), .vdd(vdd), .A(_14020_), .Y(_14021_) );
	OAI21X1 OAI21X1_5556 ( .gnd(gnd), .vdd(vdd), .A(_14021_), .B(_14016_), .C(_14825__bF_buf3), .Y(_14022_) );
	AOI21X1 AOI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_14016_), .B(_14021_), .C(_14022_), .Y(_14023_) );
	AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf2), .B(csr_9_), .Y(_14024_) );
	AOI22X1 AOI22X1_723 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_9_), .B(_14916__bF_buf3), .C(_14024_), .D(_14896__bF_buf1), .Y(_14025_) );
	OAI21X1 OAI21X1_5557 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf2), .B(_14025_), .C(_14822__bF_buf3), .Y(_14026_) );
	AOI21X1 AOI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_14017_), .C(_14789__bF_buf1), .Y(_14027_) );
	OAI21X1 OAI21X1_5558 ( .gnd(gnd), .vdd(vdd), .A(_14026_), .B(_14023_), .C(_14027_), .Y(_14028_) );
	AOI21X1 AOI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_14028_), .B(_14015_), .C(rst_bF_buf43), .Y(_13985__9_) );
	NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_14846_), .B(_14517_), .Y(_14029_) );
	NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .B(biu_ins_30_bF_buf1), .Y(_14030_) );
	OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_14029_), .B(_14030_), .Y(_14031_) );
	OAI21X1 OAI21X1_5559 ( .gnd(gnd), .vdd(vdd), .A(_14002_), .B(_14020_), .C(_14019_), .Y(_14032_) );
	INVX1 INVX1_2180 ( .gnd(gnd), .vdd(vdd), .A(_14032_), .Y(_14033_) );
	NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_14005_), .B(_14021_), .Y(_14034_) );
	OAI21X1 OAI21X1_5560 ( .gnd(gnd), .vdd(vdd), .A(_14034_), .B(_14000_), .C(_14033_), .Y(_14035_) );
	XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_14035_), .B(_14031_), .Y(_14036_) );
	AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf1), .B(csr_10_), .Y(_14037_) );
	AOI22X1 AOI22X1_724 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_10_), .B(_14916__bF_buf2), .C(_14037_), .D(_14896__bF_buf0), .Y(_14038_) );
	AOI21X1 AOI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf4), .B(_14038_), .C(_14903__bF_buf5), .Y(_14039_) );
	OAI21X1 OAI21X1_5561 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf3), .B(_14036_), .C(_14039_), .Y(_14040_) );
	AOI21X1 AOI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_10_), .C(_14789__bF_buf0), .Y(_14041_) );
	OAI21X1 OAI21X1_5562 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_10_), .B(_14324__bF_buf1), .C(_14328__bF_buf5), .Y(_14042_) );
	AOI21X1 AOI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_14040_), .B(_14041_), .C(_14042_), .Y(_13985__10_) );
	OAI21X1 OAI21X1_5563 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf0), .B(_14323__bF_buf0), .C(addr_csr_11_), .Y(_14043_) );
	INVX1 INVX1_2181 ( .gnd(gnd), .vdd(vdd), .A(_14029_), .Y(_14044_) );
	INVX1 INVX1_2182 ( .gnd(gnd), .vdd(vdd), .A(_14035_), .Y(_14045_) );
	OAI21X1 OAI21X1_5564 ( .gnd(gnd), .vdd(vdd), .A(_14030_), .B(_14045_), .C(_14044_), .Y(_14046_) );
	NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_14847_), .B(_14543_), .Y(_14047_) );
	NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_11_), .B(biu_ins_31_bF_buf6), .Y(_14048_) );
	NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_14048_), .B(_14047_), .Y(_14049_) );
	OAI21X1 OAI21X1_5565 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_14046_), .C(_14825__bF_buf1), .Y(_14050_) );
	AOI21X1 AOI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_14046_), .B(_14049_), .C(_14050_), .Y(_14051_) );
	AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf0), .B(csr_11_), .Y(_14052_) );
	AOI22X1 AOI22X1_725 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_11_), .B(_14916__bF_buf1), .C(_14052_), .D(_14896__bF_buf4), .Y(_14053_) );
	OAI21X1 OAI21X1_5566 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf0), .B(_14053_), .C(_14822__bF_buf2), .Y(_14054_) );
	AOI21X1 AOI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14847_), .C(_14789__bF_buf4), .Y(_14055_) );
	OAI21X1 OAI21X1_5567 ( .gnd(gnd), .vdd(vdd), .A(_14054_), .B(_14051_), .C(_14055_), .Y(_14056_) );
	AOI21X1 AOI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_14056_), .B(_14043_), .C(rst_bF_buf42), .Y(_13985__11_) );
	INVX1 INVX1_2183 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .Y(_14057_) );
	OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_14057_), .B(_14031_), .Y(_14058_) );
	AOI21X1 AOI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_14029_), .C(_14047_), .Y(_14059_) );
	OAI21X1 OAI21X1_5568 ( .gnd(gnd), .vdd(vdd), .A(_14033_), .B(_14058_), .C(_14059_), .Y(_14060_) );
	INVX1 INVX1_2184 ( .gnd(gnd), .vdd(vdd), .A(_14060_), .Y(_14061_) );
	NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_14034_), .B(_14058_), .Y(_14062_) );
	INVX1 INVX1_2185 ( .gnd(gnd), .vdd(vdd), .A(_14062_), .Y(_14063_) );
	OAI21X1 OAI21X1_5569 ( .gnd(gnd), .vdd(vdd), .A(_14063_), .B(_14000_), .C(_14061_), .Y(_14064_) );
	XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(csr_gpr_iu_rs1_12_), .Y(_14065_) );
	XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14064_), .B(_14065_), .Y(_14066_) );
	AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf4), .B(csr_12_), .Y(_14067_) );
	AOI22X1 AOI22X1_726 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .B(_14916__bF_buf0), .C(_14067_), .D(_14896__bF_buf3), .Y(_14068_) );
	AOI21X1 AOI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf2), .B(_14068_), .C(_14903__bF_buf2), .Y(_14069_) );
	OAI21X1 OAI21X1_5570 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf1), .B(_14066_), .C(_14069_), .Y(_14070_) );
	AOI21X1 AOI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_12_), .C(_14789__bF_buf3), .Y(_14071_) );
	OAI21X1 OAI21X1_5571 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_12_), .B(_14324__bF_buf0), .C(_14328__bF_buf4), .Y(_14072_) );
	AOI21X1 AOI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_14070_), .B(_14071_), .C(_14072_), .Y(_13985__12_) );
	OAI21X1 OAI21X1_5572 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf3), .B(_14323__bF_buf3), .C(addr_csr_13_bF_buf2), .Y(_14073_) );
	INVX1 INVX1_2186 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_12_), .Y(_14074_) );
	NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_14065_), .B(_14064_), .Y(_14075_) );
	OAI21X1 OAI21X1_5573 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14074_), .C(_14075_), .Y(_14076_) );
	NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(csr_gpr_iu_rs1_13_), .Y(_14077_) );
	INVX1 INVX1_2187 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .Y(_14078_) );
	NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14078_), .Y(_14079_) );
	NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_14077_), .B(_14079_), .Y(_14080_) );
	OAI21X1 OAI21X1_5574 ( .gnd(gnd), .vdd(vdd), .A(_14080_), .B(_14076_), .C(_14825__bF_buf4), .Y(_14081_) );
	AOI21X1 AOI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_14076_), .B(_14080_), .C(_14081_), .Y(_14082_) );
	AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(csr_13_), .Y(_14083_) );
	AOI22X1 AOI22X1_727 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_13_), .B(_14916__bF_buf3), .C(_14083_), .D(_14896__bF_buf2), .Y(_14084_) );
	OAI21X1 OAI21X1_5575 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf3), .B(_14084_), .C(_14822__bF_buf1), .Y(_14085_) );
	AOI21X1 AOI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_14078_), .C(_14789__bF_buf2), .Y(_14086_) );
	OAI21X1 OAI21X1_5576 ( .gnd(gnd), .vdd(vdd), .A(_14085_), .B(_14082_), .C(_14086_), .Y(_14087_) );
	AOI21X1 AOI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_14087_), .B(_14073_), .C(rst_bF_buf41), .Y(_13985__13_) );
	OAI22X1 OAI22X1_836 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14838_), .C(_14077_), .D(_14075_), .Y(_14088_) );
	XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(csr_gpr_iu_rs1_14_), .Y(_14089_) );
	XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_14088_), .B(_14089_), .Y(_14090_) );
	AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf2), .B(csr_14_), .Y(_14091_) );
	AOI22X1 AOI22X1_728 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_14_), .B(_14916__bF_buf2), .C(_14091_), .D(_14896__bF_buf1), .Y(_14092_) );
	AOI21X1 AOI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf0), .B(_14092_), .C(_14903__bF_buf5), .Y(_14093_) );
	OAI21X1 OAI21X1_5577 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .B(_14090_), .C(_14093_), .Y(_14094_) );
	AOI21X1 AOI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_14_), .C(_14789__bF_buf1), .Y(_14095_) );
	OAI21X1 OAI21X1_5578 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_14_), .B(_14324__bF_buf8), .C(_14328__bF_buf3), .Y(_14096_) );
	AOI21X1 AOI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_14094_), .B(_14095_), .C(_14096_), .Y(_13985__14_) );
	OAI21X1 OAI21X1_5579 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf2), .B(_14323__bF_buf2), .C(addr_csr_15_bF_buf3), .Y(_14097_) );
	NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_14089_), .B(_14088_), .Y(_14098_) );
	OAI21X1 OAI21X1_5580 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14836_), .C(_14098_), .Y(_14099_) );
	XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf2), .B(csr_gpr_iu_rs1_15_), .Y(_14100_) );
	OAI21X1 OAI21X1_5581 ( .gnd(gnd), .vdd(vdd), .A(_14100_), .B(_14099_), .C(_14825__bF_buf2), .Y(_14101_) );
	AOI21X1 AOI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_14099_), .B(_14100_), .C(_14101_), .Y(_14102_) );
	NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(csr_15_), .B(_14912__bF_buf1), .Y(_14103_) );
	NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_14103_), .B(_13990_), .Y(_14104_) );
	AOI21X1 AOI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_15_), .B(_14916__bF_buf1), .C(_14104_), .Y(_14105_) );
	OAI21X1 OAI21X1_5582 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf1), .B(_14105_), .C(_14822__bF_buf0), .Y(_14106_) );
	AOI21X1 AOI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14837_), .C(_14789__bF_buf0), .Y(_14107_) );
	OAI21X1 OAI21X1_5583 ( .gnd(gnd), .vdd(vdd), .A(_14106_), .B(_14102_), .C(_14107_), .Y(_14108_) );
	AOI21X1 AOI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_14108_), .B(_14097_), .C(rst_bF_buf40), .Y(_13985__15_) );
	NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_14065_), .B(_14080_), .Y(_14109_) );
	NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_14089_), .B(_14100_), .Y(_14110_) );
	NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_14110_), .B(_14109_), .Y(_14111_) );
	NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_14111_), .B(_14062_), .Y(_14112_) );
	AOI22X1 AOI22X1_729 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(_14839_), .C(_14111_), .D(_14060_), .Y(_14113_) );
	OAI21X1 OAI21X1_5584 ( .gnd(gnd), .vdd(vdd), .A(_14112_), .B(_14000_), .C(_14113_), .Y(_14114_) );
	XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(csr_gpr_iu_rs1_16_), .Y(_14115_) );
	XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_14114_), .B(_14115_), .Y(_14116_) );
	AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf0), .B(csr_16_), .Y(_14117_) );
	AOI22X1 AOI22X1_730 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_16_), .B(_14916__bF_buf0), .C(_14117_), .D(_14896__bF_buf0), .Y(_14118_) );
	AOI21X1 AOI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf4), .B(_14118_), .C(_14903__bF_buf2), .Y(_14119_) );
	OAI21X1 OAI21X1_5585 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf3), .B(_14116_), .C(_14119_), .Y(_14120_) );
	AOI21X1 AOI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_16_), .C(_14789__bF_buf4), .Y(_14121_) );
	OAI21X1 OAI21X1_5586 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_16_), .B(_14324__bF_buf7), .C(_14328__bF_buf2), .Y(_14122_) );
	AOI21X1 AOI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_14120_), .B(_14121_), .C(_14122_), .Y(_13985__16_) );
	OAI21X1 OAI21X1_5587 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf1), .B(_14323__bF_buf1), .C(addr_csr_17_bF_buf3), .Y(_14123_) );
	INVX1 INVX1_2188 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_16_), .Y(_14124_) );
	NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_14115_), .B(_14114_), .Y(_14125_) );
	OAI21X1 OAI21X1_5588 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14124_), .C(_14125_), .Y(_14126_) );
	XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(csr_gpr_iu_rs1_17_), .Y(_14127_) );
	INVX1 INVX1_2189 ( .gnd(gnd), .vdd(vdd), .A(_14127_), .Y(_14128_) );
	OAI21X1 OAI21X1_5589 ( .gnd(gnd), .vdd(vdd), .A(_14128_), .B(_14126_), .C(_14825__bF_buf0), .Y(_14129_) );
	AOI21X1 AOI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_14126_), .B(_14128_), .C(_14129_), .Y(_14130_) );
	AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf4), .B(csr_17_), .Y(_14131_) );
	AOI22X1 AOI22X1_731 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_17_), .B(_14916__bF_buf3), .C(_14131_), .D(_14896__bF_buf4), .Y(_14132_) );
	OAI21X1 OAI21X1_5590 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf4), .B(_14132_), .C(_14822__bF_buf3), .Y(_14133_) );
	INVX1 INVX1_2190 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_17_), .Y(_14134_) );
	AOI21X1 AOI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_14134_), .C(_14789__bF_buf3), .Y(_14135_) );
	OAI21X1 OAI21X1_5591 ( .gnd(gnd), .vdd(vdd), .A(_14133_), .B(_14130_), .C(_14135_), .Y(_14136_) );
	AOI21X1 AOI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_14136_), .B(_14123_), .C(rst_bF_buf39), .Y(_13985__17_) );
	INVX1 INVX1_2191 ( .gnd(gnd), .vdd(vdd), .A(_14114_), .Y(_14137_) );
	NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_14115_), .B(_14128_), .Y(_14138_) );
	OAI22X1 OAI22X1_837 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14829_), .C(_14138_), .D(_14137_), .Y(_14139_) );
	XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(csr_gpr_iu_rs1_18_), .Y(_14140_) );
	XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_14139_), .B(_14140_), .Y(_14141_) );
	AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(csr_18_), .Y(_14142_) );
	AOI22X1 AOI22X1_732 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_18_), .B(_14916__bF_buf2), .C(_14142_), .D(_14896__bF_buf3), .Y(_14143_) );
	AOI21X1 AOI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf2), .B(_14143_), .C(_14903__bF_buf5), .Y(_14144_) );
	OAI21X1 OAI21X1_5592 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf1), .B(_14141_), .C(_14144_), .Y(_14145_) );
	AOI21X1 AOI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_18_), .C(_14789__bF_buf2), .Y(_14146_) );
	OAI21X1 OAI21X1_5593 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_18_), .B(_14324__bF_buf6), .C(_14328__bF_buf1), .Y(_14147_) );
	AOI21X1 AOI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_14145_), .B(_14146_), .C(_14147_), .Y(_13985__18_) );
	OAI21X1 OAI21X1_5594 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf0), .B(_14323__bF_buf0), .C(addr_csr_19_bF_buf0), .Y(_14148_) );
	NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14139_), .Y(_14149_) );
	OAI21X1 OAI21X1_5595 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14827_), .C(_14149_), .Y(_14150_) );
	XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(csr_gpr_iu_rs1_19_), .Y(_14151_) );
	INVX1 INVX1_2192 ( .gnd(gnd), .vdd(vdd), .A(_14151_), .Y(_14152_) );
	OAI21X1 OAI21X1_5596 ( .gnd(gnd), .vdd(vdd), .A(_14152_), .B(_14150_), .C(_14825__bF_buf3), .Y(_14153_) );
	AOI21X1 AOI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_14150_), .B(_14152_), .C(_14153_), .Y(_14154_) );
	NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(csr_19_), .B(_14912__bF_buf2), .Y(_14155_) );
	NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_14155_), .B(_13990_), .Y(_14156_) );
	AOI21X1 AOI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_19_), .B(_14916__bF_buf1), .C(_14156_), .Y(_14157_) );
	OAI21X1 OAI21X1_5597 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf2), .B(_14157_), .C(_14822__bF_buf2), .Y(_14158_) );
	AOI21X1 AOI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14828_), .C(_14789__bF_buf1), .Y(_14159_) );
	OAI21X1 OAI21X1_5598 ( .gnd(gnd), .vdd(vdd), .A(_14158_), .B(_14154_), .C(_14159_), .Y(_14160_) );
	AOI21X1 AOI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_14160_), .B(_14148_), .C(rst_bF_buf38), .Y(_13985__19_) );
	NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14831_), .Y(_14161_) );
	NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14152_), .Y(_14162_) );
	NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_14138_), .B(_14162_), .Y(_14163_) );
	AOI21X1 AOI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_14114_), .B(_14163_), .C(_14161_), .Y(_14164_) );
	XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(csr_gpr_iu_rs1_20_), .Y(_14165_) );
	XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_14164_), .B(_14165_), .Y(_14166_) );
	AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf1), .B(csr_20_), .Y(_14167_) );
	AOI22X1 AOI22X1_733 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_20_), .B(_14916__bF_buf0), .C(_14167_), .D(_14896__bF_buf2), .Y(_14168_) );
	AOI21X1 AOI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf0), .B(_14168_), .C(_14903__bF_buf2), .Y(_14169_) );
	OAI21X1 OAI21X1_5599 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .B(_14166_), .C(_14169_), .Y(_14170_) );
	AOI21X1 AOI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_20_), .C(_14789__bF_buf0), .Y(_14171_) );
	OAI21X1 OAI21X1_5600 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_20_), .B(_14324__bF_buf5), .C(_14328__bF_buf0), .Y(_14172_) );
	AOI21X1 AOI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_14170_), .B(_14171_), .C(_14172_), .Y(_13985__20_) );
	OAI21X1 OAI21X1_5601 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf3), .B(_14323__bF_buf3), .C(addr_csr_21_bF_buf1), .Y(_14173_) );
	NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf2), .B(csr_gpr_iu_rs1_20_), .Y(_14174_) );
	INVX1 INVX1_2193 ( .gnd(gnd), .vdd(vdd), .A(_14165_), .Y(_14175_) );
	OAI21X1 OAI21X1_5602 ( .gnd(gnd), .vdd(vdd), .A(_14175_), .B(_14164_), .C(_14174_), .Y(_14176_) );
	XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(csr_gpr_iu_rs1_21_), .Y(_14177_) );
	AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_14176_), .B(_14177_), .Y(_14178_) );
	OAI21X1 OAI21X1_5603 ( .gnd(gnd), .vdd(vdd), .A(_14177_), .B(_14176_), .C(_14825__bF_buf1), .Y(_14179_) );
	OAI21X1 OAI21X1_5604 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_csrrs), .B(csr_gpr_iu_csrrw), .C(csr_gpr_iu_rs1_21_), .Y(_14180_) );
	NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(csr_21_), .B(_14912__bF_buf0), .Y(_14181_) );
	OAI21X1 OAI21X1_5605 ( .gnd(gnd), .vdd(vdd), .A(_14181_), .B(_13990_), .C(_14180_), .Y(_14182_) );
	AOI21X1 AOI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf4), .B(_14182_), .C(_14903__bF_buf0), .Y(_14183_) );
	OAI21X1 OAI21X1_5606 ( .gnd(gnd), .vdd(vdd), .A(_14178_), .B(_14179_), .C(_14183_), .Y(_14184_) );
	AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_14184_), .B(_14324__bF_buf4), .Y(_14185_) );
	OAI21X1 OAI21X1_5607 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_21_), .B(_14822__bF_buf1), .C(_14185_), .Y(_14186_) );
	AOI21X1 AOI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_14186_), .B(_14173_), .C(rst_bF_buf37), .Y(_13985__21_) );
	NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_14165_), .B(_14177_), .Y(_14187_) );
	OAI22X1 OAI22X1_838 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14832_), .C(_14187_), .D(_14164_), .Y(_14188_) );
	OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(csr_gpr_iu_rs1_22_), .Y(_14189_) );
	NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(csr_gpr_iu_rs1_22_), .Y(_14190_) );
	NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_14190_), .B(_14189_), .Y(_14191_) );
	XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_14188_), .B(_14191_), .Y(_14192_) );
	AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf4), .B(csr_22_), .Y(_14193_) );
	AOI22X1 AOI22X1_734 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_22_), .B(_14916__bF_buf3), .C(_14193_), .D(_14896__bF_buf1), .Y(_14194_) );
	AOI21X1 AOI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf3), .B(_14194_), .C(_14903__bF_buf5), .Y(_14195_) );
	OAI21X1 OAI21X1_5608 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf2), .B(_14192_), .C(_14195_), .Y(_14196_) );
	AOI21X1 AOI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_22_), .C(_14789__bF_buf4), .Y(_14197_) );
	OAI21X1 OAI21X1_5609 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_22_), .B(_14324__bF_buf3), .C(_14328__bF_buf5), .Y(_14198_) );
	AOI21X1 AOI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_14196_), .B(_14197_), .C(_14198_), .Y(_13985__22_) );
	OAI21X1 OAI21X1_5610 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf2), .B(_14323__bF_buf2), .C(addr_csr_23_bF_buf3), .Y(_14199_) );
	NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(_14189_), .B(_14190_), .C(_14188_), .Y(_14200_) );
	NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_14190_), .B(_14200_), .Y(_14201_) );
	XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(csr_gpr_iu_rs1_23_), .Y(_14202_) );
	INVX1 INVX1_2194 ( .gnd(gnd), .vdd(vdd), .A(_14202_), .Y(_14203_) );
	OAI21X1 OAI21X1_5611 ( .gnd(gnd), .vdd(vdd), .A(_14203_), .B(_14201_), .C(_14825__bF_buf0), .Y(_14204_) );
	AOI21X1 AOI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_14201_), .B(_14203_), .C(_14204_), .Y(_14205_) );
	AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(csr_23_), .Y(_14206_) );
	AOI22X1 AOI22X1_735 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_23_), .B(_14916__bF_buf2), .C(_14206_), .D(_14896__bF_buf0), .Y(_14207_) );
	OAI21X1 OAI21X1_5612 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf4), .B(_14207_), .C(_14822__bF_buf0), .Y(_14208_) );
	INVX1 INVX1_2195 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_23_), .Y(_14209_) );
	AOI21X1 AOI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14209_), .C(_14789__bF_buf3), .Y(_14210_) );
	OAI21X1 OAI21X1_5613 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_14205_), .C(_14210_), .Y(_14211_) );
	AOI21X1 AOI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_14211_), .B(_14199_), .C(rst_bF_buf36), .Y(_13985__23_) );
	NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_14191_), .B(_14187_), .Y(_14212_) );
	AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_14212_), .B(_14203_), .Y(_14213_) );
	NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_14163_), .B(_14213_), .Y(_14214_) );
	INVX1 INVX1_2196 ( .gnd(gnd), .vdd(vdd), .A(_14214_), .Y(_14215_) );
	AOI22X1 AOI22X1_736 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(_14834_), .C(_14161_), .D(_14213_), .Y(_14216_) );
	INVX1 INVX1_2197 ( .gnd(gnd), .vdd(vdd), .A(_14216_), .Y(_14217_) );
	AOI21X1 AOI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_14114_), .B(_14215_), .C(_14217_), .Y(_14218_) );
	INVX1 INVX1_2198 ( .gnd(gnd), .vdd(vdd), .A(_14218_), .Y(_14219_) );
	XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(csr_gpr_iu_rs1_24_), .Y(_14220_) );
	NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_14220_), .B(_14219_), .Y(_14221_) );
	INVX1 INVX1_2199 ( .gnd(gnd), .vdd(vdd), .A(_14221_), .Y(_14222_) );
	NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_14220_), .B(_14219_), .Y(_14223_) );
	OAI21X1 OAI21X1_5614 ( .gnd(gnd), .vdd(vdd), .A(_14223_), .B(_14222_), .C(_14825__bF_buf3), .Y(_14224_) );
	AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf2), .B(csr_24_), .Y(_14225_) );
	AOI22X1 AOI22X1_737 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_24_), .B(_14916__bF_buf1), .C(_14225_), .D(_14896__bF_buf4), .Y(_14226_) );
	AOI21X1 AOI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf1), .B(_14226_), .C(_14903__bF_buf2), .Y(_14227_) );
	NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_14227_), .B(_14224_), .Y(_14228_) );
	AOI21X1 AOI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_24_), .C(_14789__bF_buf2), .Y(_14229_) );
	OAI21X1 OAI21X1_5615 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_24_), .B(_14324__bF_buf2), .C(_14328__bF_buf4), .Y(_14230_) );
	AOI21X1 AOI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_14228_), .B(_14229_), .C(_14230_), .Y(_13985__24_) );
	OAI21X1 OAI21X1_5616 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf1), .B(_14323__bF_buf1), .C(addr_csr_25_bF_buf1), .Y(_14231_) );
	OAI21X1 OAI21X1_5617 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14840_), .C(_14221_), .Y(_14232_) );
	XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf2), .B(csr_gpr_iu_rs1_25_), .Y(_14233_) );
	AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_14232_), .B(_14233_), .Y(_14234_) );
	OAI21X1 OAI21X1_5618 ( .gnd(gnd), .vdd(vdd), .A(_14233_), .B(_14232_), .C(_14825__bF_buf2), .Y(_14235_) );
	NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(csr_25_), .B(_14912__bF_buf1), .Y(_14236_) );
	OAI22X1 OAI22X1_839 ( .gnd(gnd), .vdd(vdd), .A(_14841_), .B(_14893_), .C(_14236_), .D(_13990_), .Y(_14237_) );
	AOI21X1 AOI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf0), .B(_14237_), .C(_14903__bF_buf0), .Y(_14238_) );
	OAI21X1 OAI21X1_5619 ( .gnd(gnd), .vdd(vdd), .A(_14234_), .B(_14235_), .C(_14238_), .Y(_14239_) );
	AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_14239_), .B(_14324__bF_buf1), .Y(_14240_) );
	OAI21X1 OAI21X1_5620 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_25_), .B(_14822__bF_buf3), .C(_14240_), .Y(_14241_) );
	AOI21X1 AOI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_14241_), .B(_14231_), .C(rst_bF_buf35), .Y(_13985__25_) );
	NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_14840_), .B(_14841_), .Y(_14242_) );
	NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_14220_), .B(_14233_), .Y(_14243_) );
	INVX1 INVX1_2200 ( .gnd(gnd), .vdd(vdd), .A(_14243_), .Y(_14244_) );
	AOI22X1 AOI22X1_738 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(_14242_), .C(_14244_), .D(_14219_), .Y(_14245_) );
	OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(csr_gpr_iu_rs1_26_), .Y(_14246_) );
	NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(csr_gpr_iu_rs1_26_), .Y(_14247_) );
	AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_14246_), .B(_14247_), .Y(_14248_) );
	XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_14245_), .B(_14248_), .Y(_14249_) );
	AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf0), .B(csr_26_), .Y(_14250_) );
	AOI22X1 AOI22X1_739 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_26_), .B(_14916__bF_buf0), .C(_14250_), .D(_14896__bF_buf3), .Y(_14251_) );
	AOI21X1 AOI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .B(_14251_), .C(_14903__bF_buf5), .Y(_14252_) );
	OAI21X1 OAI21X1_5621 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf4), .B(_14249_), .C(_14252_), .Y(_14253_) );
	AOI21X1 AOI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_26_), .C(_14789__bF_buf1), .Y(_14254_) );
	OAI21X1 OAI21X1_5622 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_26_), .B(_14324__bF_buf0), .C(_14328__bF_buf3), .Y(_14255_) );
	AOI21X1 AOI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_14253_), .B(_14254_), .C(_14255_), .Y(_13985__26_) );
	OAI21X1 OAI21X1_5623 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf0), .B(_14323__bF_buf0), .C(addr_csr_27_bF_buf2), .Y(_14256_) );
	INVX1 INVX1_2201 ( .gnd(gnd), .vdd(vdd), .A(_14248_), .Y(_14257_) );
	OAI21X1 OAI21X1_5624 ( .gnd(gnd), .vdd(vdd), .A(_14257_), .B(_14245_), .C(_14247_), .Y(_14258_) );
	XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(csr_gpr_iu_rs1_27_), .Y(_14259_) );
	INVX1 INVX1_2202 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .Y(_14260_) );
	OAI21X1 OAI21X1_5625 ( .gnd(gnd), .vdd(vdd), .A(_14260_), .B(_14258_), .C(_14825__bF_buf1), .Y(_14261_) );
	AOI21X1 AOI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .B(_14260_), .C(_14261_), .Y(_14262_) );
	AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf4), .B(csr_27_), .Y(_14263_) );
	AOI22X1 AOI22X1_740 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_27_), .B(_14916__bF_buf3), .C(_14263_), .D(_14896__bF_buf2), .Y(_14264_) );
	OAI21X1 OAI21X1_5626 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf0), .B(_14264_), .C(_14822__bF_buf2), .Y(_14265_) );
	INVX1 INVX1_2203 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_27_), .Y(_14266_) );
	AOI21X1 AOI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_14266_), .C(_14789__bF_buf0), .Y(_14267_) );
	OAI21X1 OAI21X1_5627 ( .gnd(gnd), .vdd(vdd), .A(_14265_), .B(_14262_), .C(_14267_), .Y(_14268_) );
	AOI21X1 AOI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14256_), .C(rst_bF_buf34), .Y(_13985__27_) );
	NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .B(_14257_), .Y(_14269_) );
	NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_14244_), .B(_14269_), .Y(_14270_) );
	NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf4), .B(_14843_), .Y(_14271_) );
	OAI21X1 OAI21X1_5628 ( .gnd(gnd), .vdd(vdd), .A(_14270_), .B(_14218_), .C(_14271_), .Y(_14272_) );
	XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf3), .B(csr_gpr_iu_rs1_28_), .Y(_14273_) );
	INVX1 INVX1_2204 ( .gnd(gnd), .vdd(vdd), .A(_14273_), .Y(_14274_) );
	XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_14272_), .B(_14274_), .Y(_14275_) );
	AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf3), .B(csr_28_), .Y(_14276_) );
	AOI22X1 AOI22X1_741 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_28_), .B(_14916__bF_buf2), .C(_14276_), .D(_14896__bF_buf1), .Y(_14277_) );
	AOI21X1 AOI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf3), .B(_14277_), .C(_14903__bF_buf2), .Y(_14278_) );
	OAI21X1 OAI21X1_5629 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf2), .B(_14275_), .C(_14278_), .Y(_14279_) );
	AOI21X1 AOI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(csr_gpr_iu_rs1_28_), .C(_14789__bF_buf4), .Y(_14280_) );
	OAI21X1 OAI21X1_5630 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_28_), .B(_14324__bF_buf8), .C(_14328__bF_buf2), .Y(_14281_) );
	AOI21X1 AOI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_14279_), .B(_14280_), .C(_14281_), .Y(_13985__28_) );
	OAI21X1 OAI21X1_5631 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf3), .B(_14323__bF_buf3), .C(addr_csr_29_bF_buf1), .Y(_14282_) );
	INVX1 INVX1_2205 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_28_), .Y(_14283_) );
	NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_14273_), .B(_14272_), .Y(_14284_) );
	OAI21X1 OAI21X1_5632 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14283_), .C(_14284_), .Y(_14285_) );
	XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf2), .B(csr_gpr_iu_rs1_29_), .Y(_14286_) );
	INVX1 INVX1_2206 ( .gnd(gnd), .vdd(vdd), .A(_14286_), .Y(_14287_) );
	OAI21X1 OAI21X1_5633 ( .gnd(gnd), .vdd(vdd), .A(_14287_), .B(_14285_), .C(_14825__bF_buf4), .Y(_14288_) );
	AOI21X1 AOI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_14285_), .B(_14287_), .C(_14288_), .Y(_14289_) );
	AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf2), .B(csr_29_), .Y(_14290_) );
	AOI22X1 AOI22X1_742 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_29_), .B(_14916__bF_buf1), .C(_14290_), .D(_14896__bF_buf0), .Y(_14291_) );
	OAI21X1 OAI21X1_5634 ( .gnd(gnd), .vdd(vdd), .A(_14825__bF_buf3), .B(_14291_), .C(_14822__bF_buf1), .Y(_14292_) );
	INVX1 INVX1_2207 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_29_), .Y(_14293_) );
	AOI21X1 AOI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_14293_), .C(_14789__bF_buf3), .Y(_14294_) );
	OAI21X1 OAI21X1_5635 ( .gnd(gnd), .vdd(vdd), .A(_14292_), .B(_14289_), .C(_14294_), .Y(_14295_) );
	AOI21X1 AOI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_14295_), .B(_14282_), .C(rst_bF_buf33), .Y(_13985__29_) );
	INVX1 INVX1_2208 ( .gnd(gnd), .vdd(vdd), .A(_14860_), .Y(_14296_) );
	NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_14286_), .B(_14274_), .Y(_14297_) );
	AOI22X1 AOI22X1_743 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf1), .B(_14296_), .C(_14297_), .D(_14272_), .Y(_14298_) );
	OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf0), .B(csr_gpr_iu_rs1_30_), .Y(_14299_) );
	NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf6), .B(csr_gpr_iu_rs1_30_), .Y(_14300_) );
	NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14299_), .Y(_14301_) );
	XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14298_), .B(_14301_), .Y(_14302_) );
	AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_14912__bF_buf1), .B(csr_30_), .Y(_14303_) );
	AOI22X1 AOI22X1_744 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_30_), .B(_14916__bF_buf0), .C(_14303_), .D(_14896__bF_buf4), .Y(_14304_) );
	AOI21X1 AOI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf1), .B(_14304_), .C(_14903__bF_buf5), .Y(_14305_) );
	OAI21X1 OAI21X1_5636 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf0), .B(_14302_), .C(_14305_), .Y(_14306_) );
	AOI21X1 AOI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(csr_gpr_iu_rs1_30_), .C(_14789__bF_buf2), .Y(_14307_) );
	OAI21X1 OAI21X1_5637 ( .gnd(gnd), .vdd(vdd), .A(addr_csr_30_), .B(_14324__bF_buf7), .C(_14328__bF_buf1), .Y(_14308_) );
	AOI21X1 AOI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_14306_), .B(_14307_), .C(_14308_), .Y(_13985__30_) );
	OAI21X1 OAI21X1_5638 ( .gnd(gnd), .vdd(vdd), .A(_14321__bF_buf2), .B(_14323__bF_buf2), .C(addr_csr_31_bF_buf3), .Y(_14309_) );
	OAI21X1 OAI21X1_5639 ( .gnd(gnd), .vdd(vdd), .A(_14301_), .B(_14298_), .C(_14300_), .Y(_14310_) );
	XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(biu_ins_31_bF_buf5), .B(csr_gpr_iu_rs1_31_), .Y(_14311_) );
	AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_14310_), .B(_14311_), .Y(_14312_) );
	OAI21X1 OAI21X1_5640 ( .gnd(gnd), .vdd(vdd), .A(_14311_), .B(_14310_), .C(_14825__bF_buf2), .Y(_14313_) );
	INVX1 INVX1_2209 ( .gnd(gnd), .vdd(vdd), .A(csr_gpr_iu_rs1_31_), .Y(_14314_) );
	NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(csr_31_), .B(_14912__bF_buf0), .Y(_14315_) );
	OAI22X1 OAI22X1_840 ( .gnd(gnd), .vdd(vdd), .A(_14314_), .B(_14893_), .C(_14315_), .D(_13990_), .Y(_14316_) );
	AOI21X1 AOI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_14824__bF_buf5), .B(_14316_), .C(_14903__bF_buf3), .Y(_14317_) );
	OAI21X1 OAI21X1_5641 ( .gnd(gnd), .vdd(vdd), .A(_14312_), .B(_14313_), .C(_14317_), .Y(_14318_) );
	OAI21X1 OAI21X1_5642 ( .gnd(gnd), .vdd(vdd), .A(_14816_), .B(_14821_), .C(_14314_), .Y(_14319_) );
	NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(_14324__bF_buf6), .B(_14319_), .C(_14318_), .Y(_14320_) );
	AOI21X1 AOI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14309_), .C(rst_bF_buf32), .Y(_13985__31_) );
	DFFPOSX1 DFFPOSX1_1980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_13985__0_), .Q(addr_csr_0_) );
	DFFPOSX1 DFFPOSX1_1981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_13985__1_), .Q(addr_csr_1_) );
	DFFPOSX1 DFFPOSX1_1982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_13985__2_), .Q(addr_csr_2_) );
	DFFPOSX1 DFFPOSX1_1983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_13985__3_), .Q(addr_csr_3_) );
	DFFPOSX1 DFFPOSX1_1984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_13985__4_), .Q(addr_csr_4_) );
	DFFPOSX1 DFFPOSX1_1985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_13985__5_), .Q(addr_csr_5_) );
	DFFPOSX1 DFFPOSX1_1986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_13985__6_), .Q(addr_csr_6_) );
	DFFPOSX1 DFFPOSX1_1987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_13985__7_), .Q(addr_csr_7_) );
	DFFPOSX1 DFFPOSX1_1988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_13985__8_), .Q(addr_csr_8_) );
	DFFPOSX1 DFFPOSX1_1989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_13985__9_), .Q(addr_csr_9_) );
	DFFPOSX1 DFFPOSX1_1990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_13985__10_), .Q(addr_csr_10_) );
	DFFPOSX1 DFFPOSX1_1991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_13985__11_), .Q(addr_csr_11_) );
	DFFPOSX1 DFFPOSX1_1992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_13985__12_), .Q(addr_csr_12_) );
	DFFPOSX1 DFFPOSX1_1993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_13985__13_), .Q(addr_csr_13_) );
	DFFPOSX1 DFFPOSX1_1994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_13985__14_), .Q(addr_csr_14_) );
	DFFPOSX1 DFFPOSX1_1995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_13985__15_), .Q(addr_csr_15_) );
	DFFPOSX1 DFFPOSX1_1996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_13985__16_), .Q(addr_csr_16_) );
	DFFPOSX1 DFFPOSX1_1997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_13985__17_), .Q(addr_csr_17_) );
	DFFPOSX1 DFFPOSX1_1998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_13985__18_), .Q(addr_csr_18_) );
	DFFPOSX1 DFFPOSX1_1999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_13985__19_), .Q(addr_csr_19_) );
	DFFPOSX1 DFFPOSX1_2000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_13985__20_), .Q(addr_csr_20_) );
	DFFPOSX1 DFFPOSX1_2001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_13985__21_), .Q(addr_csr_21_) );
	DFFPOSX1 DFFPOSX1_2002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_13985__22_), .Q(addr_csr_22_) );
	DFFPOSX1 DFFPOSX1_2003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_13985__23_), .Q(addr_csr_23_) );
	DFFPOSX1 DFFPOSX1_2004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_13985__24_), .Q(addr_csr_24_) );
	DFFPOSX1 DFFPOSX1_2005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_13985__25_), .Q(addr_csr_25_) );
	DFFPOSX1 DFFPOSX1_2006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_13985__26_), .Q(addr_csr_26_) );
	DFFPOSX1 DFFPOSX1_2007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_13985__27_), .Q(addr_csr_27_) );
	DFFPOSX1 DFFPOSX1_2008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_13985__28_), .Q(addr_csr_28_) );
	DFFPOSX1 DFFPOSX1_2009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_13985__29_), .Q(addr_csr_29_) );
	DFFPOSX1 DFFPOSX1_2010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_13985__30_), .Q(addr_csr_30_) );
	DFFPOSX1 DFFPOSX1_2011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_13985__31_), .Q(addr_csr_31_) );
	DFFPOSX1 DFFPOSX1_2012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_13986__0_), .Q(csr_gpr_iu_csr_pc_next_0_) );
	DFFPOSX1 DFFPOSX1_2013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_13986__1_), .Q(csr_gpr_iu_csr_pc_next_1_) );
	DFFPOSX1 DFFPOSX1_2014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_13986__2_), .Q(csr_gpr_iu_csr_pc_next_2_) );
	DFFPOSX1 DFFPOSX1_2015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_13986__3_), .Q(csr_gpr_iu_csr_pc_next_3_) );
	DFFPOSX1 DFFPOSX1_2016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_13986__4_), .Q(csr_gpr_iu_csr_pc_next_4_) );
	DFFPOSX1 DFFPOSX1_2017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_13986__5_), .Q(csr_gpr_iu_csr_pc_next_5_) );
	DFFPOSX1 DFFPOSX1_2018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_13986__6_), .Q(csr_gpr_iu_csr_pc_next_6_) );
	DFFPOSX1 DFFPOSX1_2019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_13986__7_), .Q(csr_gpr_iu_csr_pc_next_7_) );
	DFFPOSX1 DFFPOSX1_2020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_13986__8_), .Q(csr_gpr_iu_csr_pc_next_8_) );
	DFFPOSX1 DFFPOSX1_2021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_13986__9_), .Q(csr_gpr_iu_csr_pc_next_9_) );
	DFFPOSX1 DFFPOSX1_2022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_13986__10_), .Q(csr_gpr_iu_csr_pc_next_10_) );
	DFFPOSX1 DFFPOSX1_2023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_13986__11_), .Q(csr_gpr_iu_csr_pc_next_11_) );
	DFFPOSX1 DFFPOSX1_2024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_13986__12_), .Q(csr_gpr_iu_csr_pc_next_12_) );
	DFFPOSX1 DFFPOSX1_2025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_13986__13_), .Q(csr_gpr_iu_csr_pc_next_13_) );
	DFFPOSX1 DFFPOSX1_2026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_13986__14_), .Q(csr_gpr_iu_csr_pc_next_14_) );
	DFFPOSX1 DFFPOSX1_2027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_13986__15_), .Q(csr_gpr_iu_csr_pc_next_15_) );
	DFFPOSX1 DFFPOSX1_2028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_13986__16_), .Q(csr_gpr_iu_csr_pc_next_16_) );
	DFFPOSX1 DFFPOSX1_2029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_13986__17_), .Q(csr_gpr_iu_csr_pc_next_17_) );
	DFFPOSX1 DFFPOSX1_2030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_13986__18_), .Q(csr_gpr_iu_csr_pc_next_18_) );
	DFFPOSX1 DFFPOSX1_2031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_13986__19_), .Q(csr_gpr_iu_csr_pc_next_19_) );
	DFFPOSX1 DFFPOSX1_2032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_13986__20_), .Q(csr_gpr_iu_csr_pc_next_20_) );
	DFFPOSX1 DFFPOSX1_2033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_13986__21_), .Q(csr_gpr_iu_csr_pc_next_21_) );
	DFFPOSX1 DFFPOSX1_2034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_13986__22_), .Q(csr_gpr_iu_csr_pc_next_22_) );
	DFFPOSX1 DFFPOSX1_2035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_13986__23_), .Q(csr_gpr_iu_csr_pc_next_23_) );
	DFFPOSX1 DFFPOSX1_2036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_13986__24_), .Q(csr_gpr_iu_csr_pc_next_24_) );
	DFFPOSX1 DFFPOSX1_2037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_13986__25_), .Q(csr_gpr_iu_csr_pc_next_25_) );
	DFFPOSX1 DFFPOSX1_2038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_13986__26_), .Q(csr_gpr_iu_csr_pc_next_26_) );
	DFFPOSX1 DFFPOSX1_2039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_13986__27_), .Q(csr_gpr_iu_csr_pc_next_27_) );
	DFFPOSX1 DFFPOSX1_2040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_13986__28_), .Q(csr_gpr_iu_csr_pc_next_28_) );
	DFFPOSX1 DFFPOSX1_2041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_13986__29_), .Q(csr_gpr_iu_csr_pc_next_29_) );
	DFFPOSX1 DFFPOSX1_2042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_13986__30_), .Q(csr_gpr_iu_csr_pc_next_30_) );
	DFFPOSX1 DFFPOSX1_2043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_13986__31_), .Q(csr_gpr_iu_csr_pc_next_31_) );
endmodule
