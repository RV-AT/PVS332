library verilog;
use verilog.vl_types.all;
entity prv332sv0_tb is
end prv332sv0_tb;
