library verilog;
use verilog.vl_types.all;
entity BUS_TB is
end BUS_TB;
